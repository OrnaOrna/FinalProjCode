`define W11_1 64'b1111100001111100001111100001111110001111110001111110001111110001
`define W11_2 64'b0111001010001011110001000010101000110001100101000110000001100011
`define W11_3 64'b1111111110111010110101001000000010010110111001010000010100001000
`define W11_4 64'b1100100000010110100001110010101110010100111010111000000001110001
`define W11_5 64'b0111111101000111000010111110111100100100011010110011110100111001
`define W11_6 64'b0111100000000110111000011111000000111010101100010101110010111111
`define W11_7 64'b1111001010111001111000111011110111110001001001111010101000011101
`define W11_8 64'b0100100000100100100110100000011001010100001010101100101011111101
`define W11_9 64'b1001100001001100001001100001001100001001000001000000001000000001
`define W11_10 64'b0011101001100111101101100110100110010101011101000111100100101111
`define W11_11 64'b0000000111110011011111010000111100010111001101100101100001110001
`define W11_12 64'b1100100001011110110100010011101001110100110111111110110101010100
`define W11_13 64'b0001100001111110000001110111000101101010001000110000000110011001
`define W11_14 64'b1000000111011000010111001111010011101101000010011101101111101001
`define W11_15 64'b0100100000100100000110100001000010110100010110101000010010100111
`define W11_16 64'b1011101000011101000011111100001101010101110010111110001001011100
`define W11_17 64'b0101110011111100100111000010101010001001001001010110010110111101
`define W11_18 64'b0110000011101001000110000110010100110100000001001000111011100101
`define W11_19 64'b1110000010100010000011111101110100110111000101001111001110101100
`define W11_20 64'b0100001111100001000101001000100111111111111100111100110101011110
`define W11_21 64'b0010100000010100110110111001110111010110100111101011101011101101
`define W11_22 64'b1101110000001011001101111111001010110110110101011100010000010100
`define W11_23 64'b1010100010101011111011110001001000100001111011101110010000100100
`define W11_24 64'b1100001110110101010010110010111001100011101010111011101101010100
`define W11_25 64'b1111001101010110001000001000101010001110001110001010010011100010
`define W11_26 64'b0101001011010010000101010110111000101000011001001010111000101010
`define W11_27 64'b1110100100110011011000000110111111101010010100100101100000010111
`define W11_28 64'b1101001001000000001011110101111100010101001001101011100000110001
`define W11_29 64'b0110100100010100001100111011011100011111000001001110111111100101
`define W11_30 64'b0011010111111100000000110011101010110101011010100010000101101110
`define W11_31 64'b0111001111101011111100111011101101100001100001111110000000010000
`define W11_32 64'b1011010111101110010111101101100100001000011110100110010110010010
`define W11_33 64'b1001101010000000010110011100110110110010000001001011111100000101
`define W11_34 64'b0100010100010011111001010001000100101011101001010110011100000001
`define W11_35 64'b0001101011011010101010110100101011011001110111110011000010111000
`define W11_36 64'b1001011110010010111101111000001101010101110010101000110100001010
`define W11_37 64'b1110001111101101001111011111010001101011110101111110011001000111
`define W11_38 64'b1100010111111000100000001011000001011010011111101111111100100110
`define W11_39 64'b0110001100110111001101100001000010000000100101101000101001100000
`define W11_40 64'b0001011100101011000100100110011111110110000001100000001001101000
`define W11_41 64'b0110000011110111000110001101110011111100101001111110101000110001
`define W11_42 64'b0111010000100000010000001001011010000011010001001110010011001010
`define W11_43 64'b0001010111110110000010001010010100100000001111100011000010011100
`define W11_44 64'b1010100001010101010110011111111011110111000001000010101011101111
`define W11_45 64'b1001010110001010101010010100000110010100110011100101001100100000
`define W11_46 64'b0010100000010100010001011011001011111110010111000110000101010011
`define W11_47 64'b1111010000101001001111010101101001000010000111000000011111011111
`define W11_48 64'b1110000001101010111100010111000000101001100111110111110110100100
`define W11_49 64'b0111010111100101011001000000001001011100000001000001000010110000
`define W11_50 64'b0001011111111001010000011101100000100110111100100111001110001011
`define W11_51 64'b1001001011100011001111000110101110110111101101010110010001110100
`define W11_52 64'b1100100000000011010010100001100110110110011011001001010110111111
`define W11_53 64'b0100100011010100010100101111100111110110001100101011100001100100
`define W11_54 64'b0001001001111100111010011011011000000111011010111100110010101111
`define W11_55 64'b1111010100011101101100010011100000001011001011110101111100011110
`define W11_56 64'b1001011100101110000001100110011101100110011001001000000100011000
`define W11_57 64'b1010001101110000000011110111011011010111110010001000101111101110
`define W11_58 64'b1101101001101111110011101100011010010011110001010010101110011100
`define W11_59 64'b0110100100001110010101100000100110101111011100100101010111101101
`define W11_60 64'b1100100010011101001010101111100001111110000011111101111111101000
`define W11_61 64'b1110100110100111100011110011100011101111000011011111011010010101
`define W11_62 64'b0010001101101000000011001001111111111110000001001111000011001100
`define W11_63 64'b0101101010001110110011011010111111000011101010100101000010111110
`define W11_64 64'b0100100000110100110100101100100100111110101110001111110010110001
`define W11_65 64'b1000011001101101101101010010001100111011101001000001011000100000
`define W11_66 64'b0110111110100100111111111100111100011101110000101101110100001010
`define W11_67 64'b0000011000100100001111010111010010111010011010001111110100001001
`define W11_68 64'b1100000111011101001111001110001110100101100001100100001110101111
`define W11_69 64'b0010011101111011110101100100011110000101010001000100001001101101
`define W11_70 64'b1110111110101010001111111101100101011011100000011011011011101011
`define W11_71 64'b1010011110010011011111110011011100100101000011100010111101100101
`define W11_72 64'b0100000101111101010100100011010011001101000001000110100111100000
`define W11_73 64'b0111000110011101011100001100110100111010001111000011000001000101
`define W11_74 64'b1110011000111101000001010010101101101011010111000001111001111100
`define W11_75 64'b0110011000001010100011011011110110010100000100001101010001111011
`define W11_76 64'b1011111110110100101010110001010110101100010000010010110101000100
`define W11_77 64'b1011100110011100001110001101010000101010111000010001101001001011
`define W11_78 64'b0011111100010100101001010001001011000100001000110100100111010010
`define W11_79 64'b0011100101110100111011111111101110001010110010110011011011110101
`define W11_80 64'b1111000111110011101100000111010100011100011000011110101101101100
`define W11_81 64'b1001011000100110001101100110000001010100111011100111110110001101
`define W11_82 64'b0010000000100011001110110011010001111001001100101011000001011101
`define W11_83 64'b1010000001010101001011010100010001000111010010000001101000000010
`define W11_84 64'b0001011011010000001000001000011011101010001000101111011101100100
`define W11_85 64'b0100000010100100101000101100101100001000100001101100001000010010
`define W11_86 64'b1000100001000000111001101000000101011010100011111001001111001010
`define W11_87 64'b0000100011001000100011100011000100011010010010111011100111110101
`define W11_88 64'b1100000000101100010010100011101101001000010000100010100011100101
`define W11_89 64'b0001001111010011101100001000001101011101010100010000101111001000
`define W11_90 64'b1001001100001111010010110110011001000110001111000010011100011101
`define W11_91 64'b0010000110101101011100110110110011010101011011100100111010101001
`define W11_92 64'b0111010110110100110101010101001010001010000100101111011100000001
`define W11_93 64'b1001110011100111001001110010010000010100101001000100111001100101
`define W11_94 64'b1111010101111011010101000111111111011001001001001110100101110101
`define W11_95 64'b1010000110110110011100101011010011010010011110011010010101011101
`define W11_96 64'b0001110010111011110100110101001010001111110110100111111000111111
`define W11_97 64'b1010010101000000011101010100010100101110000001000010001100010100
`define W11_98 64'b0010010100110100001110000010111110000011100001101010011111101111
`define W11_99 64'b0101111111000100100110100010010111011100110010010011011101010001
`define W11_100 64'b1010001110111111001000001010011000000001010001110000101100101000
`define W11_101 64'b1101111101101001111001010100111111000101100101001110110000101010
`define W11_102 64'b1011010010111001010100011100011000100101101110101011111011111010
`define W11_103 64'b0010001101101110110111110001001111100100110001011000111110001100
`define W11_104 64'b0011010001001101000011010001100000001000100111010001111110110101
`define W11_105 64'b1110100001001011110110110101011100100111101101101001111100100101
`define W11_106 64'b0110100001110101000001011011000101010001111110100101110111001100
`define W11_107 64'b0001011011101010001110100111010000101110010111000101011101101000
`define W11_108 64'b1001011001010100111001000111101011011000011011100000001100000001
`define W11_109 64'b0111011001010111110100011010101001010011111100101110010010010101
`define W11_110 64'b0011111001110011110010110010001001000001111100111010000110001101
`define W11_111 64'b1011111001111011001000111110110010000001000000011100001101110010
`define W11_112 64'b1111011001011111101110010001001010010011100000001111000010100010
`define W11_113 64'b0011111110010110000101111001100000000111011011011111111000101011
`define W11_114 64'b1010011100111100100100000000010001001110000110010110001101000111
`define W11_115 64'b1000100111101001111111111100000101111001000010110111110010100110
`define W11_116 64'b1011111110011011010101000010111110101000110111111000111011110110
`define W11_117 64'b1100010011101100010000101101100110000010011100101010100110111001
`define W11_118 64'b0010011111101101100001101101100110001011101000101010010100100101
`define W11_119 64'b0100010000100101101111100101000110010010000001000001110101011011
`define W11_120 64'b0000100100110001111000001011101110011011001110010001110111100011
`define W11_121 64'b0100000110000001000010010010010100100001010110101100001101101011
`define W11_122 64'b1101011110010000011101110100111000100110011011100111001011110110
`define W11_123 64'b0100001000100011100000101101111011001010110001101110011010100000
`define W11_124 64'b0011101011011101101111011010101011101001100010001100100111011011
`define W11_125 64'b1100000110010101000100111010000001010010100111001001011010111101
`define W11_126 64'b1011101001011111011001010111101100011010011000100110010001110101
`define W11_127 64'b1100001011110110110110101001101001111011100000000111001010110111
`define W11_128 64'b0101011111000101111110000010010101101111111010011000100000001111
`define W11_129 64'b0000100111111100000101010101110101100111001100010111110010101100
`define W11_130 64'b1000100101101011111010111001101011100001111001010010000000000001
`define W11_131 64'b1101011110011010101010100100000000110101111111100110100010010001
`define W11_132 64'b0101011100100110110101000010110001100100011111010011010010011001
`define W11_133 64'b1000011110100011110111101000101111110001110010010110000011010001
`define W11_134 64'b0010101111001100101100110001000100000001101001101010100000001000
`define W11_135 64'b1010101111110000011001100111110100001110010100001101111100101100
`define W11_136 64'b0000011100011000011101111110000011110111010010101110101100001110
`define W11_137 64'b0110111101001001111000000011101011100010000010000010100011111001
`define W11_138 64'b1101010110100010001101001111001010101000101101101010000111100011
`define W11_139 64'b1110111111101100011000010001000010111111111010011110010011011001
`define W11_140 64'b1001000111011100110011000110000000110001100101111101100001101111
`define W11_141 64'b1111010011101010110110100111011110110001000100011111100001110011
`define W11_142 64'b0111010010111011101101001011001000000011000001000101101100111100
`define W11_143 64'b0101010111001001111010101101100011000101000110010000001000011100
`define W11_144 64'b0001000110100110000000111101101100001001001010010010111000000001
`define W11_145 64'b0011100101101011001101101011111100111100100000001100110100001000
`define W11_146 64'b1110010000100001111111010001000010100100101010001101001100010100
`define W11_147 64'b0011111001110100001100000110010111000001000101000000001001000000
`define W11_148 64'b0111011110000111000001101000100011011001011010101111010010111111
`define W11_149 64'b1011100111100101101111001001011000001010001111011000011011111001
`define W11_150 64'b1111011100001001001101011000110001111100111110100000000101011101
`define W11_151 64'b0110010010010110110011101011100101110110100101010100010100111000
`define W11_152 64'b1011111011000100111101000010100000010011110011010111011111101011
`define W11_153 64'b0010010111011000001000000010110110111001111000000110001110110000
`define W11_154 64'b1111110100110111001000100000001000011010101100100001000000011001
`define W11_155 64'b0111110101000000101001111110001111010100011100000000110000010100
`define W11_156 64'b1010100111101101101110111110111100000100001100100110101010101100
`define W11_157 64'b0010100101010000100001011011010100111011100000010010111010001000
`define W11_158 64'b1010010111001100001110110111101110100011011101101010101110010100
`define W11_159 64'b0001001010110111110011110011000101010100010010110111010000101011
`define W11_160 64'b1001001010111101001101111011111100001000000110110000011101001001
`define W11_161 64'b0110010101100001010000111111010111111011010110011011001111110010
`define W11_162 64'b1001100100010001110001001111101110111100101010001010000000000001
`define W11_163 64'b1000110001000000100000011101111101001000101110101001111010010001
`define W11_164 64'b0000110001100101111101110011001110011010101010110101111101111001
`define W11_165 64'b1100001101110100100111100110001100001000000001001000000001110110
`define W11_166 64'b0001100111101110110000100000111011011101001110011001000101110000
`define W11_167 64'b1110010111111011001000001000000000000011110100010111111010011010
`define W11_168 64'b0100001101011101101010111100000010011001010101101100000100010010
`define W11_169 64'b0001001001010100100110010100010001001000010100001101000001100110
`define W11_170 64'b1001001001101111101001101110100011001101101100001010010000001110
`define W11_171 64'b1101100011000101100111110000001010110111011001000001000000010001
`define W11_172 64'b1001111101101010010110010111101000010111100000000110010000001101
`define W11_173 64'b1011000101011000001110000000111101110111000101000001010101100110
`define W11_174 64'b0101100001101100111110001110010011101010010011100010111011101011
`define W11_175 64'b0011000111110001111011101100101001101101100011111110110001101010
`define W11_176 64'b0001111111110010001111101001000110010010100110110011001110011110
`define W11_177 64'b1001001110101011001100110001000000110100111011001010000110110010
`define W11_178 64'b1010101101100010101000011100001001111001110010101000001100011101
`define W11_179 64'b0010101111101011100100101110011101010111000001111010101001110011
`define W11_180 64'b0101011100001100010110101111000010011011001110101101010011100000
`define W11_181 64'b1101101010110001000100111011100101010010000101000000001000110010
`define W11_182 64'b0001001100010111100111101101011101100110100101000001011000010101
`define W11_183 64'b0101101000010011000010111110110110100110111100101010101100101101
`define W11_184 64'b1101011111100111011001001011011101011010000101011010011100000011
`define W11_185 64'b0010011110011010000100010110110100110011000011101111111010001010
`define W11_186 64'b1011111011100010111011101110000100000001011000011111101100001000
`define W11_187 64'b0010110001110011100001110010100011000000001101111000111010110101
`define W11_188 64'b0000100100010000011011110111111011001110100101010111010011100110
`define W11_189 64'b0011111010110010111000100100011010011011111011000100111000101100
`define W11_190 64'b1000100111111110111010100101100101011101000110001100000111001011
`define W11_191 64'b1010110010111010000000101011001101011010000011110000011100101101
`define W11_192 64'b1010011101110100001100111111011010000101101111011111011110111110
`define W11_193 64'b0101101010100110010111011010110100010010110111101010010101100011
`define W11_194 64'b1101101010101011100111001000010100100001100000001000101110101100
`define W11_195 64'b1110000101011011010111110110101000111011001011001000000010000110
`define W11_196 64'b1010111101000000101000010010110001110100000010101101111010000000
`define W11_197 64'b1011100010011100001000000010100001111010011100001010110010110111
`define W11_198 64'b0110000100100011001001101101011000001000110010101110001100101000
`define W11_199 64'b0010111110010111111101110101111000100110101000100011110110101110
`define W11_200 64'b0011100001001011010110011000000001110001101011101110000010011010
`define W11_201 64'b0101001111001100110001100111101010011110010001101000111011001111
`define W11_202 64'b0000011100001000100010110100100110010011001101000011111110101010
`define W11_203 64'b1100010000000100101110111101101010001100101111100110110101110001
`define W11_204 64'b0100010000010111110011011001101100010110101110001011111011110010
`define W11_205 64'b1001010100011110011010001010001110010010010011111101000000010111
`define W11_206 64'b1101001100011110011100110011111010000110000001000101100000001000
`define W11_207 64'b0001010101001001100010111110001010011101000011011000001111010000
`define W11_208 64'b1000011110001001011011011000110110001100101001011110100110111110
`define W11_209 64'b0111000111000110100100010101010000111011000001001111001111011001
`define W11_210 64'b1000001100001001000111110010111100101011000101110110100001011011
`define W11_211 64'b1000111101111011100010110001111100100000001111010001110000010000
`define W11_212 64'b1111000101010101011011100011101000110000000000111000001110000111
`define W11_213 64'b0000111101001001010110100111000101111000111010010110001101100000
`define W11_214 64'b0000001100110100110000011100111001110000110000000001100000100100
`define W11_215 64'b0101110001010001010000000011011100001001110010001111100001010111
`define W11_216 64'b1101110000011110010011101000010111110011001111101111100111111000
`define W11_217 64'b0011111101000000010010001010010001100000000011010000001001000001
`define W11_218 64'b0010100101011001001000000111111011101111000100011101110001111010
`define W11_219 64'b0110101010011111010000001110101100001000110110111010010000001001
`define W11_220 64'b0111001001111001000110010001000011100101111001101011100111010101
`define W11_221 64'b1010100111011010001100011101000111011000001111000100100000101110
`define W11_222 64'b1110101010011100011110000101110010100111010100010000111111100010
`define W11_223 64'b1111001011010011101000011100110100100000110010111101111111011010
`define W11_224 64'b1011111111111100000110100111100100100101010100101001011010101010
`define W11_225 64'b0010100101111011001010111011100101001010111001101010000001000011
`define W11_226 64'b0111011100100011101101000110101110001110011101011001100110001101
`define W11_227 64'b1111011101001010110010100010010111101000100001100111010110110110
`define W11_228 64'b1010100101101111110101011111011100000101111010001110010111101011
`define W11_229 64'b1001100111100001100100000000100000010000100010100010010010110000
`define W11_230 64'b1111110111101101111110111100000000010011001100111011010001011011
`define W11_231 64'b0111110101111001111110001111001110000010110000001010111101101010
`define W11_232 64'b0001100101101100010001110110111111110110101101001100100010011000
`define W11_233 64'b0100000101010111001010001100011011011000000101010100111100000111
`define W11_234 64'b1011100110101101110010010001000110010111000001001101001011010100
`define W11_235 64'b1111011101100000111101101101111000010000010110101100010101110110
`define W11_236 64'b1100000101101100001111010010000101101001011001011111101100110000
`define W11_237 64'b0111011111011000100101110011010111011010010100100111000101000001
`define W11_238 64'b0000110010011111001100100110111011010110100010011010001111011110
`define W11_239 64'b0011100101100010110111110100001101100100101101011001000100010100
`define W11_240 64'b1000110000101000111001101000010110100110001110001001101101100101
