`define L1 64'b1000000001000000001000000001000000001000000001000000001000000001
`define L2 64'b1000000011000000101000001111000010001000110011001010101011111111
`define L3 64'b1000000000010010011001010001000110111010100100111010010100001010
`define L4 64'b1000000011010100100011110010111000000110011001001100000010111110
`define L5 64'b1000000011010100100001010000100001000011110010011001110010101100
`define L6 64'b1000000011110010001001111101001011100111010110010010111111100010
`define L7 64'b1000000000110000000010101110100000100111100100110001101011101110
`define L8 64'b1000000001010000001000100110100000111001001001011101001000001110
`define L9 64'b1000000001110100110111010001101010110101010110010101110010100100
`define L10 64'b1000000011010100001011011011101010110010111011001111101011011000
`define L11 64'b1000000000000100101100111010110100001100111110001101101000010100
`define L12 64'b1000000001101000101001100001010001001001101011011010111110001101
`define L13 64'b1000000011101000010001100011110010110111100110110011000100111011
`define L14 64'b1000000011100100010000011001011101011010101001100100010010011100
`define L15 64'b1000000001100000001010000001111011101001001111101111000100110100
`define L16 64'b1000000011001100111111000000011111110110011110101110000010011001
`define L17 64'b1000000000000100110001010001101101010011101110000101110101000111
`define L18 64'b1000000011100000101010001101011001110001001010010100101111111001
`define L19 64'b1000000011001100111100111111010001110010010101110011110010110110
`define L20 64'b1000000001101100010001111001111100010001000001000010011000101110
`define L21 64'b1000000011011000001011111100011011010100111011110111001001100001
`define L22 64'b1000000010111000001101111011101010100111000101010000010001011011
`define L23 64'b1000000000100100010110010110000100001111110011001100011001001110
`define L24 64'b1000000000000100010001011101110000111010101010010001010010110110
`define L25 64'b1000000001011000110010011111001010111001110000111100110011101101
`define L26 64'b1000000000111000101100010010011001111100111100010011101010011111
`define L27 64'b1000000011100000101010001101011001101111110101110001110101100111
`define L28 64'b1000000000000100010101001001100101110110101100101110000000000111
`define L29 64'b1000000000000100011111000010100011111001010011111010011101011000
`define L30 64'b1000000001100000001010000001111010010111101111101110111110011100
