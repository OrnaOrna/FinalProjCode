// Parameters used by the RAMBAM module with d=4 and P,Q chosen as per the original paper
`define P 9'b110101001
`define Q 5'b10001
`define PQ 13'b1101100111001
`define d 4
`define W 144'b010111000000111111000000100111000000001010100000100010010000001001010000011001010000101111010000101011110000100011000000001011100000011010010000
`define w 12'b101001000000
`define pow1 144'b100000000000001000000000000010000000000000100000000000001000000000000010110110011100001101100111101110001011100110110000001001101100000010011011
`define pow2 144'b100000000000000010000000000000001000110110011100101110001011001001101100101101110100011001111001000111010100011011010011111100100101101000010011
`define pow4 144'b100000000000101110001011000111010100111111101001101011111101111000010111110000100110010000101110010011010001101000100000001010100000101101000111
`define L 64'b1000000000010010011001010001000110111010100100111010010100001010
`define L_inv 64'b1000000010100010010111011101010010010101000110111001010011000100
`define modPmat 32'b11010100011010100011010111001110
`define mulL2 144'b000100100000000010010000000001001000000000100100000000010010000000001001110110011000011011001100001101100110000110110011110101000101101100111110