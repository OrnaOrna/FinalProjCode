`define P1 9'b110110001
`define P2 9'b101110001
`define P3 9'b110101001
`define P4 9'b101101001
`define P5 9'b100111001
`define P6 9'b111111001
`define P7 9'b101100101
`define P8 9'b111110101
`define P9 9'b110001101
`define P10 9'b101001101
`define P11 9'b100101101
`define P12 9'b100011101
`define P13 9'b111011101
`define P14 9'b110111101
`define P15 9'b111000011
`define P16 9'b110100011
`define P17 9'b101100011
`define P18 9'b111110011
`define P19 9'b110001011
`define P20 9'b100101011
`define P21 9'b100011011
`define P22 9'b101111011
`define P23 9'b110000111
`define P24 9'b111100111
`define P25 9'b111010111
`define P26 9'b101110111
`define P27 9'b111001111
`define P28 9'b110011111
`define P29 9'b101011111
`define P30 9'b100111111
