`define W21_1 64'b1100110001100110001100111001100101111000100010000100010010010110
`define W21_2 64'b0011101010000110001011000000001111110001010011101010101001110111
`define W21_3 64'b1000101101110001100000100000000011111101000111001111110100000000
`define W21_4 64'b1011100110000010111100010101010110111010010101101000000101101101
`define W21_5 64'b0010101101101111100001001101010001010000000101001110110001000011
`define W21_6 64'b0110110000000000110010100011001001010101100001110010101000101010
`define W21_7 64'b1101111111100000111001011110000000011001101101001011000111000110
`define W21_8 64'b1110011010101100010010100111111001101000101011001101001000101110
`define W21_9 64'b0001110000001110000001110000001100011101000100100001010100001010
`define W21_10 64'b1100100010110011000000000101110000000000001001010000000011000001
`define W21_11 64'b1101110010000001001010100000011111101001000111110010110111011100
`define W21_12 64'b1110111110010011101110010100101100101001111100100010101000110100
`define W21_13 64'b1011110000011010011000011101110101000101000110011100010000111110
`define W21_14 64'b0111110010010100010011011101100010101000000011010111110011101001
`define W21_15 64'b0100111010000110010111100111111011010010001100000001000000000000
`define W21_16 64'b1001101100011100010111011010000101111011000101010011101010111101
`define W21_17 64'b0111101111100110000110111010011111111010001001101001101000100110
`define W21_18 64'b0011110000100001101010011111100111111001000110011011000010001000
`define W21_19 64'b0101111100000011010111110101110010000001111000010000001100101100
`define W21_20 64'b0000110010101101000001011010110111110010001100011001000010100100
`define W21_21 64'b1110101111001001000000000000000001100001110010011001110101100110
`define W21_22 64'b0010010000100100001100011011111001011110000000100100100101011110
`define W21_23 64'b0010101111101011000000101110011000001101001001011100111000000001
`define W21_24 64'b0010011101001100101011111100101111011101100111100110101100000000
`define W21_25 64'b1101010110101100010110011101010101101111010100110000101001111001
`define W21_26 64'b1111100101100000010111100100101111000111111011000111111011010010
`define W21_27 64'b0000000010110100111000100111001100011010101000101001110101011010
`define W21_28 64'b0011000011101000000000001110011101111111001000101000010110100111
`define W21_29 64'b0101110100001001111000000001011100010111010110011010111000011010
`define W21_30 64'b1101001000001000100111111011010111111001010011000100110000000001
`define W21_31 64'b0000100010001011001010001100001000010001101100101010001110100011
`define W21_32 64'b1111110000000000100100110010110011110100100000101011011111110100
`define W21_33 64'b0111110111000111110000000001100100000100011110101010001111011001
`define W21_34 64'b0100011010110100000000010010001011010001010100101111001011110010
`define W21_35 64'b1100101010100010110110110001101100000000011010000101000001111001
`define W21_36 64'b0001011111001110100111010000000010001111100010101101110000011001
`define W21_37 64'b0011011111111001011011000111000111101011011100010000000010110000
`define W21_38 64'b1100110101101101000000001011011111010101110110100010011101000101
`define W21_39 64'b1111100111100101011011010001000011110101111000110001000011101001
`define W21_40 64'b0001110010010111010110010000001000011100110100001100110000101110
`define W21_41 64'b1111010011111100011110111011011110000111000010000001110001110011
`define W21_42 64'b1011100110101011000000001101100111110100011111111110011011110100
`define W21_43 64'b1010110000001011001000001010010000011010000100101000110010100100
`define W21_44 64'b0101010101010101101011101000001000111001011010001110101011111011
`define W21_45 64'b0101000100010101111111100010011001100010000000001110110011011111
`define W21_46 64'b1001010101011110010110001010100001010100111110100000101000111101
`define W21_47 64'b0001100001101001110111101101101111111000011011001010111101010010
`define W21_48 64'b0100000101011110110100010100000101111111100011110101010101010101
`define W21_49 64'b1011000101010010101000010101001001010110010100101010011100010000
`define W21_50 64'b0100111111010101111101101001101000100011101010011100100000000000
`define W21_51 64'b0001001100010010000000011011111010101101011010011100101000001111
`define W21_52 64'b1011110001001010000000001011110010010111110101101111011000100010
`define W21_53 64'b1110100111100110010100111000001101110010001110011100011111101001
`define W21_54 64'b0011001100111011100110100011110011110101110011100011001111000001
`define W21_55 64'b1001000101101001001010000011011101101001100100101100110011001100
`define W21_56 64'b1100010101101110111011011111101000011001010001100011000111011100
`define W21_57 64'b0000110010000101110111111001011010100110101101011001011010011010
`define W21_58 64'b1111111111010000101101001110100010100101101100101000101001011100
`define W21_59 64'b0011100000011100110100010110111110000011100001101100110111110000
`define W21_60 64'b1101110010101011100111100000101000001011010000101101011001001000
`define W21_61 64'b0001101000011010100001111011110000010011110101011111010001111010
`define W21_62 64'b0010110010110000100010111111011001101110010101010100011001111001
`define W21_63 64'b1101111101000110101110100111000111101101101010110010001101000110
`define W21_64 64'b0101111101100101000000000111100010011011101100001110111101000010
`define W21_65 64'b1001111110001101000110000001001000000110101111100010000100000110
`define W21_66 64'b0001001011101111000110010011011100100101001101111100011000001011
`define W21_67 64'b0111000110001110000000000010100101010000101110101000111010010011
`define W21_68 64'b0001111101101110010111100010111100011111101100101101111100011100
`define W21_69 64'b1001110011100001010100011010011101111101111101101111011001111011
`define W21_70 64'b1011010010101011100010001000010111110101001111000010111010010111
`define W21_71 64'b1101001111000101110011110001110000101101111101000111100001101110
`define W21_72 64'b1001011111000101001000001011001100100000111110000001100110101110
`define W21_73 64'b1010101101110110100011010011100011111011110010010101101000000000
`define W21_74 64'b0000011100100111001111000100001101100100010110100011110001100100
`define W21_75 64'b1000100101001011110000100111101111000011110101111110011100100101
`define W21_76 64'b1101111010011011101101000000010110100100101100010101000011001011
`define W21_77 64'b1101110001001010101011001011011111011100101101001010111101101000
`define W21_78 64'b0101011011001110110011001011110110000101100001010010010100011101
`define W21_79 64'b1000110100011111001101001011011010011101101110011001001011001111
`define W21_80 64'b0110110101010010100001000011111100101011101100111001000010100111
`define W21_81 64'b1111001111001001100000110011010110011010101011110001100100111010
`define W21_82 64'b0000000011111100011100010110101010100000001011011000010010100000
`define W21_83 64'b0010000001000001011000100010110101101111001000110001101100101101
`define W21_84 64'b1101001111100010100100000101001011110101001101111011000000110111
`define W21_85 64'b0101100100110111010010100111010101101110111001001110110011010011
`define W21_86 64'b1000001100001000000001011000101110010100100001101000011011011100
`define W21_87 64'b0101110111010101010010000001001001111011010010000000011110001111
`define W21_88 64'b0000011111100010110011111110010010001001011010101010010111001000
`define W21_89 64'b1001101000000110110010101100011000000011010111110000011001010011
`define W21_90 64'b0100000001001110000100100110010001010010000000000000000100101010
`define W21_91 64'b0101101001100011111011011110110100001001000010010100010101000101
`define W21_92 64'b1001010000010111100101001100000110010101010101000011010100000000
`define W21_93 64'b1110110000101111110000111001001100011100110111110000000000110100
`define W21_94 64'b0110111110000100100001001111000010111110110100000010000111101010
`define W21_95 64'b0010000101110000100010001010100100000011001011001000010111011010
`define W21_96 64'b1011100101100111000010001010001001010001000100111000011111011110
`define W21_97 64'b0111011100110100011001010010010100100001010000000010001000010010
`define W21_98 64'b0110010110011010100000100010011111010001111101100101101000010001
`define W21_99 64'b1100110110100011111100110001001010110001111010101111100001110111
`define W21_100 64'b1001111100101010000000000110000011110110001010010010100100100011
`define W21_101 64'b0000000011100110100100101100111111000111111011100101111100101011
`define W21_102 64'b1001001110100111010111101000101001000101100010100100010110001010
`define W21_103 64'b1101001000010011110000100110001010100011011100101101000111111111
`define W21_104 64'b0001000000011000100111000010110100010000100110010001100000011000
`define W21_105 64'b0010010011010100100100110010000111011010011011010000010100000101
`define W21_106 64'b1000010000100101011011001100101110100111101001111011011111101110
`define W21_107 64'b0111001111110010011010011111111111111111000110101010011101101001
`define W21_108 64'b1101001101101011000101100000001100010100110001100110101100010100
`define W21_109 64'b0001000000111001110111111011101011001111010111001110000101110010
`define W21_110 64'b1010001001001001101000111011111101111010101000110000000011101011
`define W21_111 64'b1011010000000110111111000111010110110001111111111000110000000000
`define W21_112 64'b1000011011001000110010001000011000111010011101101110110100100111
`define W21_113 64'b0111010000011101101011010100001111011001011001101100010010000111
`define W21_114 64'b1010110101110101100101111101100011100010110110000101001011001100
`define W21_115 64'b1101100001111111000000001010111110101111011110010111100001111000
`define W21_116 64'b0110011111110111000111000101100010101111000011110001001101110100
`define W21_117 64'b0011001000110101000101000010000101110110000100110011001010001101
`define W21_118 64'b1000100001001010101001100100101011001000111011011110011000000000
`define W21_119 64'b0110010111011111100110100100000111000100100000011010000101000001
`define W21_120 64'b1101101011000000001110000011110110001100010011000110101110010011
`define W21_121 64'b0101111110011110110111000000000100011100110111001110100100000000
`define W21_122 64'b0010111010000111111001001110010001010111011000110110001101011110
`define W21_123 64'b1100111011001101011000111000101100101010110000100100101001000110
`define W21_124 64'b0100011110100110000011011001110100101010001010101001110100001101
`define W21_125 64'b1001100000100100001111110100000100111111101010111010011110111100
`define W21_126 64'b0011101001110010001110100010010100100101000111110111111100001011
`define W21_127 64'b1100100011110111000000111000101011001011111101111100011010111011
`define W21_128 64'b0110100101010011010100111000101100001111000000011101011011100010
`define W21_129 64'b0101110011000010101011011010101100010111110100110011001111110001
`define W21_130 64'b0100100000000000110000111000101001000001111010001000001001000001
`define W21_131 64'b0001110110101010111001110010011111100000100101110100101010010111
`define W21_132 64'b1000011110110001010100000010001111100001100001111000011111111110
`define W21_133 64'b1011001000110011111110011100110110000110001010011100101011010000
`define W21_134 64'b0011000010110100100011001000010100101111101101001001101010101011
`define W21_135 64'b0010110111110110111000100000011011110000101001001010001010011011
`define W21_136 64'b0010111101111000100111101100100111010000101111100000000011101001
`define W21_137 64'b0001111000011011001111010010001100001001110100100011100011011011
`define W21_138 64'b0000001100000101010000101111001110100011010101100101001100000110
`define W21_139 64'b1110110101011010101001111100001101001010001011100000000000001011
`define W21_140 64'b0100011011101100000000000110111000110110101110111010010100001111
`define W21_141 64'b1000100000010011110110001001101100110111001100011111101001010000
`define W21_142 64'b0000111111001001101011010110000000000000101000101010110110011011
`define W21_143 64'b1000111011010101000001110000001001000001000110100101101100011000
`define W21_144 64'b1001111010111100010101001001111100000001001000100111100010010001
`define W21_145 64'b0001111111101101010111011101100110000100100100101000110100011111
`define W21_146 64'b1011110011010001000110010000100111011000101111000111000100000000
`define W21_147 64'b1101101111111111110110111011110010011010010100011010110010101100
`define W21_148 64'b1110000011110111111101110101111000010110011110010110111100100111
`define W21_149 64'b0101110111100000000000101101101100000000101111110001100010111101
`define W21_150 64'b1001110011000011000101100110001000101011110000001111110100010110
`define W21_151 64'b1001101011100101100110111101011011011100100100010011100101000110
`define W21_152 64'b1001100110111100101110100000000001101110011010001111011111101010
`define W21_153 64'b1100110110000101110100000100000111000100001111011001100000111101
`define W21_154 64'b1100000110110110000110101101101101100111000010100111010100010000
`define W21_155 64'b0110111110111101010110111100100110111101111111011000011101110100
`define W21_156 64'b0100110110000100100001000101111001111011100001000011011001100100
`define W21_157 64'b0000000000001111101001100010111110011010101110011011010100000000
`define W21_158 64'b1010100100100111110110111011000010101001101010011001011101110000
`define W21_159 64'b1101011000001011100000010000000001111101011001010001100011001110
`define W21_160 64'b1110101000010010010100100001001001001000111011111110101010111000
`define W21_161 64'b1011100001110101010101001111101011000100101110001010011101101010
`define W21_162 64'b0000000101011110000110001111001000011001111100111011101101010000
`define W21_163 64'b0110001001000000111011011101000010110010101000010000000011110010
`define W21_164 64'b1100100100011110111011000111111000111011011001101010100110010100
`define W21_165 64'b0011010010000010110010011111100101001111000001001011011001110111
`define W21_166 64'b0000000000000000000000000110111110111010100001110111101111011111
`define W21_167 64'b0010000000110010110101011111111011100111110101011000001000000000
`define W21_168 64'b0001001110011111110001000001010000001001000000000001001100011101
`define W21_169 64'b0000110010001010100100100010101101011000011111111001001010011110
`define W21_170 64'b0001001000010010010011001011101111010111001000000111000101001100
`define W21_171 64'b0011101001100000000000100100100010101111100001111000010100010000
`define W21_172 64'b1001101100100110101011101011000101111001111000100010011001101010
`define W21_173 64'b0011111001000001010001100000011101110111001110010001000000000000
`define W21_174 64'b1011011011101010010111001001001011101010010010101111010011010000
`define W21_175 64'b0010000001001011111011100001101010010001111101001000010111000000
`define W21_176 64'b1001101010011101001010000000001000110001000111100000001000011011
`define W21_177 64'b1110100010100011010110001100011101001011110001111001110000000000
`define W21_178 64'b1001010000101011111011000110010000110111000111001011011000100010
`define W21_179 64'b1101101010110001001011100011011101000101110110010100011000110111
`define W21_180 64'b1010110001111011010011010100010110100101000010001001101011011111
`define W21_181 64'b1001100001101001011010111111000111010000001100011101001001001000
`define W21_182 64'b1100010000111001100001000001010001101110111111101001000010111110
`define W21_183 64'b0000110001011000100000101000100101010011100001010101001111110110
`define W21_184 64'b0101011110110110000000100100000100000000111101010101001011110010
`define W21_185 64'b0100011001100000010110111000101110010110001001101110000100110001
`define W21_186 64'b0101001111001110110011100110010000110110100101001100111100000001
`define W21_187 64'b0011100011101000101101000001001101100100010001001100100001011100
`define W21_188 64'b0110100100111001001001100101000010110000100010011111100011100000
`define W21_189 64'b1011100101100001001101110011011100011010000111011011111001100001
`define W21_190 64'b0011110110011111011010000011010000011100000000001011011110110111
`define W21_191 64'b0111111001111011110111010101100111110100111100010010100100101100
`define W21_192 64'b1010110001011111001100100100101000000110000100111010110011000001
`define W21_193 64'b1001111000000000111000111111110011100110000001010101101101011110
`define W21_194 64'b0000000011101011011000100001110001011010000011010001000101000110
`define W21_195 64'b0011001110000010000001010110000111001110000000001111110110101010
`define W21_196 64'b1000111110111101001011110101110101010011111000000100111001000000
`define W21_197 64'b1000111010101000110000101110001000000110001000000111001000100000
`define W21_198 64'b0100110000001000011001010100110001001010000010001010001110001010
`define W21_199 64'b0001000101010110110011111111000010011001000010011101111011001111
`define W21_200 64'b1100101000011001101000010110000000111010100100001011100000000000
`define W21_201 64'b1000101101110111010000100101111101000010011011010001110111010100
`define W21_202 64'b0111100001101001001011001011101011100011110100110011000010110111
`define W21_203 64'b1000111001001110000010100010101100110100000101011000010010001110
`define W21_204 64'b1111001101111110011111100111100010100100000111101111010101100000
`define W21_205 64'b1011000010011010011000011100011101001000111110000010100111111011
`define W21_206 64'b1111001100000100011100000000100101010111101000000010101011111110
`define W21_207 64'b0000100110111111000000000001010011011000101000100100110110010101
`define W21_208 64'b0000011111001001010011011110110001110110010010100101010011001001
`define W21_209 64'b1110111110110101010001000110100101011010010111101010101100101101
`define W21_210 64'b0101011000101111000000000111011000000011010101100100010100110011
`define W21_211 64'b1010100100111001000011011000001110111000000000001001110110100100
`define W21_212 64'b0010101001011100101011001100111110000001111000101000000100010010
`define W21_213 64'b0001000100000011000110001111011000010001000100101110010010010100
`define W21_214 64'b1110110110011001000101100000000000101001110001000011111110000011
`define W21_215 64'b1100110100110111111010101111101000010000011000001110101100110111
`define W21_216 64'b0101010011110011010111101010110100111010111100010011000010100101
`define W21_217 64'b1001111010111111101111010000000011111101111101101111011000100011
`define W21_218 64'b1110011101001110011000100011100100000000110111100010000001011011
`define W21_219 64'b0100010010001010111110111100011000101100111000100101110100011001
`define W21_220 64'b1010101100100110110110110110111100110110111111010001000011001011
`define W21_221 64'b0011111011101000011000111000101111010110101001001111111100010111
`define W21_222 64'b1010001010011101110001011111101011111010000000000010101101101010
`define W21_223 64'b0000000011011011100000010111010011001001111101011100111101011100
`define W21_224 64'b1100011100101000100000111000001110010100011111101101010111010000
`define W21_225 64'b1110001001110010001110011010000011101001101000101001001001001001
`define W21_226 64'b1000001111111101011110111000001110011011011000110001100000010010
`define W21_227 64'b0011111101000010101101111100101010010111100111010011111100001010
`define W21_228 64'b0011000000011001110111000001010000001011110111001100100011111000
`define W21_229 64'b1010100000001000100111110001100000011001101010011011100110101000
`define W21_230 64'b0110011011000000100010101001000100010000101001100111110111000000
`define W21_231 64'b1010110101110101010011001101100001101011001001011101101001010010
`define W21_232 64'b1110001101010011011110101001110001100010111111100101001110011001
`define W21_233 64'b1001110100000000110011111100111101001011110001111100000101001011
`define W21_234 64'b1010001011010101100110111110100001001110010010100111001011010000
`define W21_235 64'b0100111110011001111011100100011000010001001100011101011000101001
`define W21_236 64'b1011100001011100010100000100110110101001001100010010000010010100
`define W21_237 64'b0110010101001010111111011100010010000100110001000100000001111001
`define W21_238 64'b1101111100101101000100111110000100000001100011001111001101010011
`define W21_239 64'b1011000111001000101100010001110110101100110010001001001101001110
`define W21_240 64'b1111011011110001000000000110111110100010111101100101001100001100
