`define W21_1 32'b10001101100100111001110000011011
`define W21_2 32'b01111001100011111111010011001001
`define W21_3 32'b11101010110010010110101100101100
`define W21_4 32'b00000000100101110001010100010110
`define W21_5 32'b10011011111100111001110111101100
`define W21_6 32'b01010110110111000001101000001010
`define W21_7 32'b00111001001100010000010100100111
`define W21_8 32'b11010111110110010011101011010101
`define W21_9 32'b10110110000000010000000001000000
`define W21_10 32'b10010110101111101001100101000010
`define W21_11 32'b11000100001000111001000101011011
`define W21_12 32'b10101000111111011101101110100010
`define W21_13 32'b01010001100010110111100001101001
`define W21_14 32'b00001000010010011000100001111001
`define W21_15 32'b11111001111000000110100010011010
`define W21_16 32'b11111100010101010010001111100100
`define W21_17 32'b10100011011001010010011000110110
`define W21_18 32'b10000100111111011110010111100100
`define W21_19 32'b01100101111101010111010000101101
`define W21_20 32'b10010101100101111110011111110001
`define W21_21 32'b11101111011001000110011001010100
`define W21_22 32'b01000101100111011010101010111001
`define W21_23 32'b11110000110110101101001011110111
`define W21_24 32'b01011000000001111111001110110111
`define W21_25 32'b10000011011010000101101011000110
`define W21_26 32'b10011100001111011001110101110001
`define W21_27 32'b00010100001111010001001001010000
`define W21_28 32'b01001000000011101111000000110011
`define W21_29 32'b01011000100111110101000010001011
`define W21_30 32'b00010001110000111011010011101000
