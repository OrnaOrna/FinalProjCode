`define W21_1 56'b10110011101011011010001000100101000010101001110110111010
`define W21_2 56'b11100011000101010110111001010011111010011011010010011010
`define W21_3 56'b11001101111011100100110000001011111111111010001101011111
`define W21_4 56'b10000011000101001001011010010101110111000010110110100110
`define W21_5 56'b01010101001111010101001100100010011010110011111111110011
`define W21_6 56'b00111100101101100111000001100000001111101000011001110101
`define W21_7 56'b00101000001000000001010000110110111010001000000111110000
`define W21_8 56'b01110101011110111001100001110111000101001101010001100100
`define W21_9 56'b01000100111100111111001010110010100000111110111100011010
`define W21_10 56'b10111000100100001011011101101100100110000001011101111100
`define W21_11 56'b10101100010010111111100100110011101000101000100010100111
`define W21_12 56'b11101001101111001001101011100011100100101001010011100000
`define W21_13 56'b11001100000101101110010111110100001101100011010010001001
`define W21_14 56'b11010011100100100101001110100010101001101011000001010110
`define W21_15 56'b10100000101110010011000111000011010101111110111110101111
`define W21_16 56'b11011100011101010000001111000100110101001100001101001100
`define W21_17 56'b00100001111001111010010010110100000000110111001111001001
`define W21_18 56'b00010010011010110111001101110010101011100000111000100000
`define W21_19 56'b11001101010111011101110010000101011100111111010110100010
`define W21_20 56'b10011110100111001110110011111010101010010011101100111110
`define W21_21 56'b01001011110000001100001011110000100000001101101101011010
`define W21_22 56'b10000000010110000110111101111100010110101110101011110001
`define W21_23 56'b11110011110110011101000111110100001001010100010010101010
`define W21_24 56'b00100010011111011000100111001101100110100000111100101001
`define W21_25 56'b00100100110011111111110101100001110100010110011111111000
`define W21_26 56'b10110000000100011011000101011101100000110111011001101011
`define W21_27 56'b11010101111111001101001110010001011100100001111011011111
`define W21_28 56'b00110101011100111000110101001110100011000101011100111111
`define W21_29 56'b10110111011100001011111101100100000011001111100000111000
`define W21_30 56'b10011111010011010011101001100110110011000101011111000101
