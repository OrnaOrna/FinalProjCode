`define w1 16'b1100011000000000
`define w2 16'b1001101110000000
`define w3 16'b1010110000000000
`define w4 16'b1011111010000000
`define w5 16'b1001110000000000
`define w6 16'b1100101100000000
`define w7 16'b1111010000000000
`define w8 16'b1011010010000000
`define w9 16'b1001111010000000
`define w10 16'b1001010100000000
`define w11 16'b1101110010000000
`define w12 16'b1011111010000000
`define w13 16'b1001110100000000
`define w14 16'b1000110010000000
`define w15 16'b1001110010000000
`define w16 16'b1101110000000000
`define w17 16'b1010010000000000
`define w18 16'b1100110000000000
`define w19 16'b1011100000000000
`define w20 16'b1010000110000000
`define w21 16'b1001010110000000
`define w22 16'b1000011100000000
`define w23 16'b1000101010000000
`define w24 16'b1011110100000000
`define w25 16'b1111000000000000
`define w26 16'b1111111100000000
`define w27 16'b1101100110000000
`define w28 16'b1000110110000000
`define w29 16'b1100110000000000
`define w30 16'b1001000100000000
`define w31 16'b1001100010000000
`define w32 16'b1010101000000000
`define w33 16'b1001110110000000
`define w34 16'b1000110010000000
`define w35 16'b1011101110000000
`define w36 16'b1101101100000000
`define w37 16'b1001111010000000
`define w38 16'b1110010000000000
`define w39 16'b1000111100000000
`define w40 16'b1001100010000000
`define w41 16'b1111100010000000
`define w42 16'b1110110000000000
`define w43 16'b1001011110000000
`define w44 16'b1101111000000000
`define w45 16'b1010001100000000
`define w46 16'b1100001110000000
`define w47 16'b1110010110000000
`define w48 16'b1010010010000000
`define w49 16'b1000101110000000
`define w50 16'b1000111000000000
`define w51 16'b1101110000000000
`define w52 16'b1100010000000000
`define w53 16'b1100000100000000
`define w54 16'b1000110010000000
`define w55 16'b1101000110000000
`define w56 16'b1011001100000000
`define w57 16'b1101110110000000
`define w58 16'b1111010000000000
`define w59 16'b1001010010000000
`define w60 16'b1000110000000000
`define w61 16'b1000010100000000
`define w62 16'b1100111110000000
`define w63 16'b1011111000000000
`define w64 16'b1011111100000000
`define w65 16'b1111000100000000
`define w66 16'b1010110010000000
`define w67 16'b1011100100000000
`define w68 16'b1000001110000000
`define w69 16'b1011000100000000
`define w70 16'b1000110000000000
`define w71 16'b1011000010000000
`define w72 16'b1010110000000000
`define w73 16'b1110010010000000
`define w74 16'b1110111100000000
`define w75 16'b1010011100000000
`define w76 16'b1111001100000000
`define w77 16'b1111011000000000
`define w78 16'b1100001010000000
`define w79 16'b1000100110000000
`define w80 16'b1100010000000000
`define w81 16'b1010011000000000
`define w82 16'b1101100100000000
`define w83 16'b1100011100000000
`define w84 16'b1101000010000000
`define w85 16'b1111010010000000
`define w86 16'b1001010100000000
`define w87 16'b1101010110000000
`define w88 16'b1100101000000000
`define w89 16'b1110101000000000
`define w90 16'b1000001100000000
`define w91 16'b1010010010000000
`define w92 16'b1100010010000000
`define w93 16'b1100001000000000
`define w94 16'b1111011100000000
`define w95 16'b1100110000000000
`define w96 16'b1111111010000000
`define w97 16'b1100001000000000
`define w98 16'b1101010100000000
`define w99 16'b1000001000000000
`define w100 16'b1110001000000000
`define w101 16'b1110101010000000
`define w102 16'b1001000000000000
`define w103 16'b1000100100000000
`define w104 16'b1110101000000000
`define w105 16'b1000011000000000
`define w106 16'b1110011000000000
`define w107 16'b1110101100000000
`define w108 16'b1110001110000000
`define w109 16'b1110001010000000
`define w110 16'b1001100110000000
`define w111 16'b1000011110000000
`define w112 16'b1100101010000000
`define w113 16'b1100111010000000
`define w114 16'b1010010100000000
`define w115 16'b1001111100000000
`define w116 16'b1100110000000000
`define w117 16'b1001111010000000
`define w118 16'b1110100000000000
`define w119 16'b1010100010000000
`define w120 16'b1000011100000000
`define w121 16'b1101011000000000
`define w122 16'b1011010100000000
`define w123 16'b1111000000000000
`define w124 16'b1011110000000000
`define w125 16'b1100001100000000
`define w126 16'b1010101000000000
`define w127 16'b1101101010000000
`define w128 16'b1100110100000000
`define w129 16'b1101000010000000
`define w130 16'b1100110100000000
`define w131 16'b1001010110000000
`define w132 16'b1001101110000000
`define w133 16'b1010111110000000
`define w134 16'b1100000110000000
`define w135 16'b1010111000000000
`define w136 16'b1110001000000000
`define w137 16'b1111101110000000
`define w138 16'b1010101110000000
`define w139 16'b1010001100000000
`define w140 16'b1110100110000000
`define w141 16'b1000100110000000
`define w142 16'b1111011110000000
`define w143 16'b1100111010000000
`define w144 16'b1101001110000000
`define w145 16'b1110001010000000
`define w146 16'b1001001110000000
`define w147 16'b1001000110000000
`define w148 16'b1101100110000000
`define w149 16'b1011010000000000
`define w150 16'b1000001110000000
`define w151 16'b1001010010000000
`define w152 16'b1101111110000000
`define w153 16'b1100111000000000
`define w154 16'b1001110010000000
`define w155 16'b1010101110000000
`define w156 16'b1001111110000000
`define w157 16'b1101001000000000
`define w158 16'b1111010100000000
`define w159 16'b1010010110000000
`define w160 16'b1111000110000000
`define w161 16'b1100010100000000
`define w162 16'b1001010000000000
`define w163 16'b1110011110000000
`define w164 16'b1100110000000000
`define w165 16'b1101001110000000
`define w166 16'b1111000010000000
`define w167 16'b1001111100000000
`define w168 16'b1100101100000000
`define w169 16'b1001010010000000
`define w170 16'b1100000000000000
`define w171 16'b1000100000000000
`define w172 16'b1001111000000000
`define w173 16'b1010000000000000
`define w174 16'b1011100010000000
`define w175 16'b1110011100000000
`define w176 16'b1000000010000000
`define w177 16'b1010111000000000
`define w178 16'b1011010010000000
`define w179 16'b1011111000000000
`define w180 16'b1110000110000000
`define w181 16'b1010110000000000
`define w182 16'b1110000010000000
`define w183 16'b1001001110000000
`define w184 16'b1101100110000000
`define w185 16'b1100101010000000
`define w186 16'b1111110000000000
`define w187 16'b1010010110000000
`define w188 16'b1011010000000000
`define w189 16'b1101001000000000
`define w190 16'b1010011000000000
`define w191 16'b1100111100000000
`define w192 16'b1110111110000000
`define w193 16'b1101011100000000
`define w194 16'b1010101110000000
`define w195 16'b1110101100000000
`define w196 16'b1001001010000000
`define w197 16'b1101100010000000
`define w198 16'b1001111000000000
`define w199 16'b1100101110000000
`define w200 16'b1110001110000000
`define w201 16'b1100100010000000
`define w202 16'b1011110000000000
`define w203 16'b1111100110000000
`define w204 16'b1011111110000000
`define w205 16'b1001110100000000
`define w206 16'b1101101010000000
`define w207 16'b1101111000000000
`define w208 16'b1001000010000000
`define w209 16'b1010101000000000
`define w210 16'b1001101000000000
`define w211 16'b1111000000000000
`define w212 16'b1001001010000000
`define w213 16'b1000001000000000
`define w214 16'b1100100100000000
`define w215 16'b1110111000000000
`define w216 16'b1001000000000000
`define w217 16'b1101011000000000
`define w218 16'b1110001100000000
`define w219 16'b1101111110000000
`define w220 16'b1001010000000000
`define w221 16'b1111101100000000
`define w222 16'b1101110100000000
`define w223 16'b1100110110000000
`define w224 16'b1101101010000000
`define w225 16'b1100001110000000
`define w226 16'b1001111100000000
`define w227 16'b1111101100000000
`define w228 16'b1000001000000000
`define w229 16'b1110010110000000
`define w230 16'b1100111000000000
`define w231 16'b1001000000000000
`define w232 16'b1011000110000000
`define w233 16'b1011000100000000
`define w234 16'b1000110010000000
`define w235 16'b1111111010000000
`define w236 16'b1001101110000000
`define w237 16'b1000011010000000
`define w238 16'b1011011100000000
`define w239 16'b1111011110000000
`define w240 16'b1000000100000000
