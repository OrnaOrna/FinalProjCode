`define W21_1 64'b1100110001100110001100111001100101111000100010000100010010010110
`define W21_2 64'b0001110000001110000001110000001100011101000100100001010100001010
`define W21_3 64'b0111101111100110000110111010011111111010001001101001101000100110
`define W21_4 64'b1101010110101100010110011101010101101111010100110000101001111001
`define W21_5 64'b0111110111000111110000000001100100000100011110101010001111011001
`define W21_6 64'b1111010011111100011110111011011110000111000010000001110001110011
`define W21_7 64'b1011000101010010101000010101001001010110010100101010011100010000
`define W21_8 64'b0000110010000101110111111001011010100110101101011001011010011010
`define W21_9 64'b1001111110001101000110000001001000000110101111100010000100000110
`define W21_10 64'b1010101101110110100011010011100011111011110010010101101000000000
`define W21_11 64'b1111001111001001100000110011010110011010101011110001100100111010
`define W21_12 64'b1001101000000110110010101100011000000011010111110000011001010011
`define W21_13 64'b0111011100110100011001010010010100100001010000000010001000010010
`define W21_14 64'b0010010011010100100100110010000111011010011011010000010100000101
`define W21_15 64'b0111010000011101101011010100001111011001011001101100010010000111
`define W21_16 64'b0101111110011110110111000000000100011100110111001110100100000000
`define W21_17 64'b0101110011000010101011011010101100010111110100110011001111110001
`define W21_18 64'b0001111000011011001111010010001100001001110100100011100011011011
`define W21_19 64'b0001111111101101010111011101100110000100100100101000110100011111
`define W21_20 64'b1100110110000101110100000100000111000100001111011001100000111101
`define W21_21 64'b1011100001110101010101001111101011000100101110001010011101101010
`define W21_22 64'b0000110010001010100100100010101101011000011111111001001010011110
`define W21_23 64'b1110100010100011010110001100011101001011110001111001110000000000
`define W21_24 64'b0100011001100000010110111000101110010110001001101110000100110001
`define W21_25 64'b1001111000000000111000111111110011100110000001010101101101011110
`define W21_26 64'b1000101101110111010000100101111101000010011011010001110111010100
`define W21_27 64'b1110111110110101010001000110100101011010010111101010101100101101
`define W21_28 64'b1001111010111111101111010000000011111101111101101111011000100011
`define W21_29 64'b1110001001110010001110011010000011101001101000101001001001001001
`define W21_30 64'b1001110100000000110011111100111101001011110001111100000101001011
