`define W21_1 24'b100101101000100010000111
`define W21_2 24'b011011101001100011100011
`define W21_3 24'b001001000000011110100101
`define W21_4 24'b101000100011010110110111
`define W21_5 24'b000101000111110000010010
`define W21_6 24'b101101010011111111111001
`define W21_7 24'b011101100111111001001010
`define W21_8 24'b101101011011101101011000
`define W21_9 24'b000010111011110010111101
`define W21_10 24'b011101110101111101111000
`define W21_11 24'b000010111110110001011110
`define W21_12 24'b011100000010010100000011
`define W21_13 24'b110101010000111111111100
`define W21_14 24'b101000101110001100100010
`define W21_15 24'b010011000101010111011101
`define W21_16 24'b011010111100001010110100
`define W21_17 24'b011100001011011011110101
`define W21_18 24'b001000000101100101000001
`define W21_19 24'b001011101011111000111111
`define W21_20 24'b111010001110101010011010
`define W21_21 24'b100110110001000000010010
`define W21_22 24'b001000111111101111001100
`define W21_23 24'b000110110011000100111001
`define W21_24 24'b100010011101011000100010
`define W21_25 24'b010011111010010010010110
`define W21_26 24'b000111101011111100011111
`define W21_27 24'b001100010001100000110111
`define W21_28 24'b011000100010010011011010
`define W21_29 24'b011001101010000101101110
`define W21_30 24'b001001011111011110000000

