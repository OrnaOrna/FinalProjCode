`define w1 14'b11000110000000
`define w2 14'b10011110100000
`define w3 14'b10100100000000
`define w4 14'b11110000000000
`define w5 14'b10011101100000
`define w6 14'b11111000100000
`define w7 14'b10001011100000
`define w8 14'b11011101100000
`define w9 14'b11110001000000
`define w10 14'b11100100100000
`define w11 14'b10100110000000
`define w12 14'b11101010000000
`define w13 14'b11000010000000
`define w14 14'b10000110000000
`define w15 14'b11001110100000
`define w16 14'b11010110000000
`define w17 14'b11010000100000
`define w18 14'b11111011100000
`define w19 14'b11100010100000
`define w20 14'b11001110000000
`define w21 14'b11000101000000
`define w22 14'b10010100100000
`define w23 14'b10101110000000
`define w24 14'b11001010100000
`define w25 14'b11010111000000
`define w26 14'b11001000100000
`define w27 14'b10101010000000
`define w28 14'b11010110000000
`define w29 14'b11000011100000
`define w30 14'b10110001000000