`define W21_1 16'b1010000010111110
`define W21_2 16'b0100000010110110
`define W21_3 16'b0001000100110010
`define W21_4 16'b1000111100011000
`define W21_5 16'b0011001101011011
`define W21_6 16'b1000101000000000
`define W21_7 16'b1110100011100000
`define W21_8 16'b0111000101111111
`define W21_9 16'b1111110001001011
`define W21_10 16'b1111100011010000
`define W21_11 16'b1011100001011111
`define W21_12 16'b1101110110001000
`define W21_13 16'b0000000011011010
`define W21_14 16'b0100101100001010
`define W21_15 16'b1110010111111100
`define W21_16 16'b1110011001001111
`define W21_17 16'b1011010101110011
`define W21_18 16'b1001101111100010
`define W21_19 16'b1011100000101000
`define W21_20 16'b0001001000010000
`define W21_21 16'b0111001111111000
`define W21_22 16'b1110111100110111
`define W21_23 16'b0100101001100000
`define W21_24 16'b1100110010010011
`define W21_25 16'b0000000011101011
`define W21_26 16'b0110110111001100
`define W21_27 16'b0111101101010010
`define W21_28 16'b0011011001110000
`define W21_29 16'b0001101011011101
`define W21_30 16'b0100110110011111
