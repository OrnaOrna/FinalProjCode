`define L1 64'b1000000001000000001000000001000000001000000001000000001000000001
`define L2 64'b1000000000100000000010000000001011011000001101101101010101011001
`define L3 64'b1000000000001000110110001101010101111010111010011100110110100011
`define L4 64'b1000000011011000011110101100110100100111001010010001011100000100
`define L5 64'b1000000010110010010111110101001001000000010110011111011100101001
`define L6 64'b1000000001111010001001110001011110110010100010011011100000110110
`define L7 64'b1000000000100111101100101011100001011111000000010101001011101001
`define L8 64'b1000000001011111010000001111011100100000101000110001000010001001
`define L9 64'b1000000011000000101000001111000010001000110011001010101011111111
`define L10 64'b1000000010100000100010001010101000111000001101101000001101000111
`define L11 64'b1000000010001000001110001000001110110010100101111111101101110101
`define L12 64'b1000000000111000101100101111101100111001110101110110100111001100
`define L13 64'b1000000010110010001110010110100101111010111101110101100000110110
`define L14 64'b1000000001111010001000011001101011000000010001111000100111010111
`define L15 64'b1000000000100001110000001000100110100000011101011111000011110111
`define L16 64'b1000000000111001011110100101100000100001111111111001101010010111
`define L17 64'b1000000000010010011001010001000110111010100100111010010100001010
`define L18 64'b1000000010111010001110010001101001111001010001111011000101001010
`define L19 64'b1000000001010001100001011010011000010010101100111101101011010101
`define L20 64'b1000000001011001010100010100111010000101000010101010011001000111
`define L21 64'b1000000000111001011110011011000101011001110101010010110110010011
`define L22 64'b1000000001111001010110010010110101010001001100000100111001000010
`define L23 64'b1000000010000101000100101101101001100101010010100001000100110000
`define L24 64'b1000000001100101101110101010010100111001010000100001101010110011
`define L25 64'b1000000011010100100011110010111000000110011001001100000010111110
`define L26 64'b1000000001111100101100111000100010010101001101110011010001100100
`define L27 64'b1000000000000110011111001010000010110011011000111000100001110001
`define L28 64'b1000000011100110110101001110111110001111011100010010111000111000
`define L29 64'b1000000011100001111001100011101011010100010000101110111100110111
`define L30 64'b1000000010010101111000010010011111100110101111100011101001100011
`define L31 64'b1000000010110011100101010011010011100001001110000010011100000101
`define L32 64'b1000000010001111000001101100000001111100000001011010000001000010
`define L33 64'b1000000011010100100001010000100001000011110010011001110010101100
`define L34 64'b1000000001111100100100010100111001100110101011000100000000111110
`define L35 64'b1000000010000110011111001111000110010001011011110100111011011000
`define L36 64'b1000000001100110110101000010000010000101001101010000100001101111
`define L37 64'b1000000010010001011001100100000011010100001100110010000001101010
`define L38 64'b1000000010000101010000111001110000011111110110000011100100110011
`define L39 64'b1000000001000011000111110011100110000110001111100111001000110101
`define L40 64'b1000000000011111100001100111001001111100011010101111000111001001
`define L41 64'b1000000011110010001001111101001011100111010110010010111111100010
`define L42 64'b1000000001011010010100110000111111110010001001010001001100100010
`define L43 64'b1000000001010011111100100001001100100111011010101101001010000101
`define L44 64'b1000000010110011010110101001001001010011111000100000111101010000
`define L45 64'b1000000001000111110011110010111010110011001000100100011001011001
`define L46 64'b1000000000100111111001110010111101000111100000110001101100100101
`define L47 64'b1000000011100111010001110001101111001111010100000010111001101010
`define L48 64'b1000000011001111101100110100011001011010100001011001001010000011
`define L49 64'b1000000000110000000010101110100000100111100100110001101011101110
`define L50 64'b1000000010011000001100000011010100001010011111101110100001001001
`define L51 64'b1000000001111000100110001100001000110000000100010011010111000011
`define L52 64'b1000000000001010001001110001101001111111011010110010010100010001
`define L53 64'b1000000001101101011110000100010110011000111011101100001001110011
`define L54 64'b1000000000100111011111110010010111101111011100111110101001111110
`define L55 64'b1000000011101111011011011000111101111000010010010100010101101011
`define L56 64'b1000000001111111111011111110101001101101110000111000111110010011
`define L57 64'b1000000001010000001000100110100000111001001001011101001000001110
`define L58 64'b1000000000011000111110001110101001010000000011110110001100010101
`define L59 64'b1000000011111000010100000110001100100010011111100110100010110111
`define L60 64'b1000000000100010001110011101001010000001101111011001001100001111
`define L61 64'b1000000010000001111100011100001011011011000101011001000100100101
`define L62 64'b1000000011110001110110111001000100011000101101111111001110111101
`define L63 64'b1000000000111001100000011001001111110001110001011100001001111110
`define L64 64'b1000000011011011000110001111001111111000000011101110101011000101
`define L65 64'b1000000001110100110111010001101010110101010110010101110010100100
`define L66 64'b1000000001111100000110111111001001111010101001000011001000111000
`define L67 64'b1000000001011010011111001011101100011011100100011111001011000010
`define L68 64'b1000000001111010011101001001001011011101101001010001101010010001
`define L69 64'b1000000010110101010110110001001101011010001110001011110010100101
`define L70 64'b1000000011011101101101010101110001011011110000100001001101111111
`define L71 64'b1000000000011011011110100011001001110100011111111001001011001100
`define L72 64'b1000000001011011010110101011110001111100110011001011101101011001
`define L73 64'b1000000011010100001011011011101010110010111011001111101011011000
`define L74 64'b1000000001011100000010111101001011100011010001110111010011101100
`define L75 64'b1000000000010010110101000000110100101101100011111011101011101010
`define L76 64'b1000000010110010010111001101101000001011000100111101001010001111
`define L77 64'b1000000000101101101100101111101001011100100000011101101000000100
`define L78 64'b1000000011101101000100101001010011010100000001000000110101000111
`define L79 64'b1000000011100011111011011010010100010010110110001001010000010011
`define L80 64'b1000000000001011111000110111010011101101111010101010010110000001
`define L81 64'b1000000000000100101100111010110100001100111110001101101000010100
`define L82 64'b1000000001000100100100110111001100000100101100011010110010101011
`define L83 64'b1000000000001100001001011100010111001100001011110110010011111101
`define L84 64'b1000000011001100100001011001101101000100100110001001001000111100
`define L85 64'b1000000010000101010001001001001010010011000101000111001100101111
`define L86 64'b1000000000100101110011000110010010000101101010111001101111111000
`define L87 64'b1000000010010011000001001010110010110011111111011010110110011000
`define L88 64'b1000000010110011000011001101101000100101001111001100010110110001
`define L89 64'b1000000001101000101001100001010001001001101011011010111110001101
`define L90 64'b1000000000111100001010011001101110011101010001000111101110110000
`define L91 64'b1000000010111010011010001101010110100110000001000001010001000100
`define L92 64'b1000000010100110010010011010111110110101101100001101110010111000
`define L93 64'b1000000001001001101101011101110000111100100010101000000100000100
`define L94 64'b1000000000101001100111010111101110111010100011011101001110001010
`define L95 64'b1000000010110101001111001000000100101001011000101001101110101101
`define L96 64'b1000000010011101101110101101001101101000101110001101010101100010
`define L97 64'b1000000011101000010001100011110010110111100110110011000100111011
`define L98 64'b1000000000010100110101111010110111001011000011000100110111010000
`define L99 64'b1000000011110010111010001000001101000110110011000011110000001100
`define L100 64'b1000000001000110101101110011000111100011110100001111010001011000
`define L101 64'b1000000011100011000101000111111111010111110010101010110110011011
`define L102 64'b1000000011001011111100101110010111101000010110001000001111001010
`define L103 64'b1000000011010111110010110100110111110010001110111110010110100010
`define L104 64'b1000000010110111111000111111010000010100101000100111111111001100
`define L105 64'b1000000011100100010000011001011101011010101001100100010010011100
`define L106 64'b1000000000101100001111111110100100010010010001100000110000110100
`define L107 64'b1000000000010010010101110011011111100100101101011100110010000111
`define L108 64'b1000000001011010101010011100100100101100111000110000010000011001
`define L109 64'b1000000001000001010110100100010010101001001101001100100110110101
`define L110 64'b1000000010101001001011000000010000111111100001111110100110100110
`define L111 64'b1000000001010111111001001100110001000001000110011001011101000110
`define L112 64'b1000000000111111000100100000110001010111100111000011011111100011
`define L113 64'b1000000001100000001010000001111011101001001111101111000100110100
`define L114 64'b1000000000101000111010011111000100010111111110011111010010100011
`define L115 64'b1000000001101100011000000010110100101000011011010001111001011101
`define L116 64'b1000000001001110110100111110010101000111010111010101111111111001
`define L117 64'b1000000011101001000101111111010001001110000101010000001101101101
`define L118 64'b1000000011010011010001110101111101101100001101001000111100010101
`define L119 64'b1000000001000111011011001000111101100000101000110010110111110101
`define L120 64'b1000000000010111010011100000001111010011111101011110010100111110
`define L121 64'b1000000011001100111111000000011111110110011110101110000010011001
`define L122 64'b1000000011111100111101101110000010111101011000011010100010100100
`define L123 64'b1000000011110110101111011010100000100001110111110101100100000101
`define L124 64'b1000000000111110110011001011010011111100000001010000011111101111
`define L125 64'b1000000000100001111111110000010010011011111011111000110101100001
`define L126 64'b1000000010111101001000010101100111111111100100110000010001111010
`define L127 64'b1000000010011011001111100010101111001100101001001011010010010011
`define L128 64'b1000000011111111100110111000110100111110100110010010101111011111
`define L129 64'b1000000000000100110001010001101101010011101110000101110101000111
`define L130 64'b1000000011010100011001111011100100000011100101000000110100111011
`define L131 64'b1000000011001100110101000010100001100111110100011011100110111000
`define L132 64'b1000000011101110000001001111100011000101010111110001101110010100
`define L133 64'b1000000011000101010100110101110111001100001110110110000000001011
`define L134 64'b1000000000000011111011100100001000000100000010111111100011010001
`define L135 64'b1000000001010011110011000110000011010100010101010010100001011111
`define L136 64'b1000000001100111000000110000110111101110010001110100001001010101
`define L137 64'b1000000011100000101010001101011001110001001010010100101111111001
`define L138 64'b1000000010101000011100010100101111000111000111000110011010111110
`define L139 64'b1000000010100100001100110100110110110101000010001000111100011100
`define L140 64'b1000000011011100111000001000010110101000100110101101011000001000
`define L141 64'b1000000001110001110001110110011010100100010000001100000110011010
`define L142 64'b1000000010110101110111000111110111100000101111101000010100100000
`define L143 64'b1000000000110011101101011000111111011100111110010111110101000000
`define L144 64'b1000000011000111101001001100000100110011001000000100110100101001
`define L145 64'b1000000011001100111100111111010001110010010101110011110010110110
`define L146 64'b1000000001110010110010100101100110000101011110111101111111111001
`define L147 64'b1000000011001010100001011101111100101110001101110010100101010111
`define L148 64'b1000000000101110101110111111010110010111101101100000010001111011
`define L149 64'b1000000010000101001011100010100110111011010001001111010101101100
`define L150 64'b1000000011110011011100100011110011001010011011000101100111111100
`define L151 64'b1000000010111011100101110000010011001100111111001001011000110111
`define L152 64'b1000000010010111110011001001011011110011111110011111010001000100
`define L153 64'b1000000001101100010001111001111100010001000001000010011000101110
`define L154 64'b1000000001100010100000111101011101001011011110001001001100000100
`define L155 64'b1000000011101110011011000011100001000111110011111001111110111111
`define L156 64'b1000000001111110111011101101010101101100110011000011100001111000
`define L157 64'b1000000000010001011000100101100110000011100101001101011111001111
`define L158 64'b1000000010000011010010111001001101111110101111110100100111111010
`define L159 64'b1000000001001011011111100100100111101110001011101101010110010100
`define L160 64'b1000000001000111000100010010011001100010111110100101100111001100
`define L161 64'b1000000011011000001011111100011011010100111011110111001001100001
`define L162 64'b1000000011010100010010100001000010010111110000100000001010111100
`define L163 64'b1000000001001010100101110000001011010011100110100011101011101111
`define L164 64'b1000000000110110110110000100110100101111101111001100011000110101
`define L165 64'b1000000011010011000110111011110100110110011000010110110011000010
`define L166 64'b1000000000011011001101100110110011011000101010110100110110011010
`define L167 64'b1000000010010111110100110011101000011011001101011011110101110100
`define L168 64'b1000000000101111110101000111001001001010011101000001000010101011
`define L169 64'b1000000010111000001101111011101010100111000101010000010001011011
`define L170 64'b1000000010010110011111011111000000001001011111001010101010011100
`define L171 64'b1000000000001001111011110000011010111000111111101111111111001011
`define L172 64'b1000000000100101100101101101000101111101110010111111000000010101
`define L173 64'b1000000001111101000010011010101011101111010110110000011011110011
`define L174 64'b1000000010100111001001011100110010010110111100111101000111101000
`define L175 64'b1000000000110111101001110000010000100101100111001100110011111110
`define L176 64'b1000000011101111101110001111111100110111111010001011101001111100
`define L177 64'b1000000000100100010110010110000100001111110011001100011001001110
`define L178 64'b1000000011001010110101010010100100011101000110000010010111001100
`define L179 64'b1000000000001110001001001101100001011001010100010110000111000001
`define L180 64'b1000000001111110000011101000001100100100000001001101100000011000
`define L181 64'b1000000001011001000011111100011011001010001100100100011100000100
`define L182 64'b1000000011010101000111010010010101111110110000011011011100110010
`define L183 64'b1000000000011101011111101011011100001110010011101000001110111100
`define L184 64'b1000000000001111110010100100011111010101101111000010100101010001
`define L185 64'b1000000000000100010001011101110000111010101010010001010010110110
`define L186 64'b1000000001100010101100111010000101001110110010011101011110101001
`define L187 64'b1000000000111010011000100100011110110011010011011010000101100111
`define L188 64'b1000000001001110000011010010001111101001101101101100110001001101
`define L189 64'b1000000011101001000001000001011001000101011001111101110000001100
`define L190 64'b1000000001000101001110100001010001100010001001000100011101010100
`define L191 64'b1000000000001101111010011100110000000100010101000001011011001001
`define L192 64'b1000000010110011010011101101011100001101000011000010001100100100
`define L193 64'b1000000001011000110010011111001010111001110000111100110011101101
`define L194 64'b1000000000010110001010110001000001110111110101000000001000110100
`define L195 64'b1000000011110001010110000000000111001001011010001111001011010100
`define L196 64'b1000000011001001101110011100110010010011001101000000010011111110
`define L197 64'b1000000010111001100100110000010000010110010001010100111101101000
`define L198 64'b1000000010010011000101100100111100101011100111010001000011000011
`define L199 64'b1000000000101011011101110000001011110001111011010110011001000101
`define L200 64'b1000000001110111111100010110011001011000111111100000000110011101
`define L201 64'b1000000000111000101100010010011001111100111100010011101010011111
`define L202 64'b1000000001111100111000101111000011101001111010101010101010010100
`define L203 64'b1000000011100010111010011010101011100101010100100111001011110001
`define L204 64'b1000000000110110001110000111101110110001100101000010011001100011
`define L205 64'b1000000010110001011111000011101011100010010111001111000011111101
`define L206 64'b1000000011101001111001010111001000101101011000110110101101011100
`define L207 64'b1000000011100101001011010110101100110110100111110010010011101010
`define L208 64'b1000000000101101001101100010010000111000111111010111101101010010
`define L209 64'b1000000011100000101010001101011001101111110101110001110101100111
`define L210 64'b1000000010101000011011110001110111011001101101000000011000111110
`define L211 64'b1000000011110100111000001011001110101000010100101101011010001000
`define L212 64'b1000000011101100000001010111101111100011100010001001000110110100
`define L213 64'b1000000011011001111011001011111100000101101000000111101111010111
`define L214 64'b1000000000000101111000111001000111110100011001110010101111000000
`define L215 64'b1000000011100011111101000010101111100000001111101011001110100000
`define L216 64'b1000000001101111110110010000011011101100110000001011111101010010
`define L217 64'b1000000000000100010101001001100101110110101100101110000000000111
`define L218 64'b1000000001010100011101101110000001101011100111111010100011101100
`define L219 64'b1000000001110110011010111010100001011111101000010100011100110011
`define L220 64'b1000000010111110000001000001110001010100001100111001100111110001
`define L221 64'b1000000000000001101011010011101110111110000001110111110110100001
`define L222 64'b1000000010101101101111100111110100000100111011000001110000100101
`define L223 64'b1000000001101011010111110100011100000001001001011100110010110010
`define L224 64'b1000000001011111000000011100110010101101111100010011101110011111
`define L225 64'b1000000000000100011111000010100011111001010011111010011101011000
`define L226 64'b1000000011001100011100110010110101100101010110001000101101011001
`define L227 64'b1000000001111100111110011010011101010101101111001011101110001101
`define L228 64'b1000000000001110110011001001100001110011001000010010110110111100
`define L229 64'b1000000011111001010101011011101100001110010110010110101000000011
`define L230 64'b1000000001100101000001000110000001111100000000110010100000100001
`define L231 64'b1000000001010101000011100110101011001100110111011001100001001111
`define L232 64'b1000000001110011011001011000101100000100100011010110000011011101
`define L233 64'b1000000001100000001010000001111010010111101111101110111110011100
`define L234 64'b1000000000101000100101111110111101101001011001111101110001110101
`define L235 64'b1000000000100100011000000001101100101000110110110001111010001011
`define L236 64'b1000000000101110111001011101001101011001100010110010000101100111
`define L237 64'b1000000001101001001011100101010111100101001000111101001110111110
`define L238 64'b1000000001011001001001001001000101100000011101010001101100100011
`define L239 64'b1000000011100101010110010010000100100100100111001001000111000011
`define L240 64'b1000000010010111011010011101110000101110110000110101010111011011
