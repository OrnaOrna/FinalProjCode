`define w1 10'b1100011000
`define w2 10'b1001111010
`define w3 10'b1010010000
`define w4 10'b1111000000
`define w5 10'b1001110110
`define w6 10'b1111100010
`define w7 10'b1000101110
`define w8 10'b1101110110
`define w9 10'b1111000100
`define w10 10'b1110010010
`define w11 10'b1010011000
`define w12 10'b1110101000
`define w13 10'b1100001000
`define w14 10'b1000011000
`define w15 10'b1100111010
`define w16 10'b1101011000
`define w17 10'b1101000010
`define w18 10'b1111101110
`define w19 10'b1110001010
`define w20 10'b1100111000
`define w21 10'b1100010100
`define w22 10'b1001010010
`define w23 10'b1010111000
`define w24 10'b1100101010
`define w25 10'b1101011100
`define w26 10'b1100100010
`define w27 10'b1010101000
`define w28 10'b1101011000
`define w29 10'b1100001110
`define w30 10'b1011000100