`define Linv1 64'b1000000001000000001000000001000000001000000001000000001000000001
`define Linv2 64'b1000000001011111010000001111011100100000101000110001000010001001
`define Linv3 64'b1000000010110010010111110101001001000000010110011111011100101001
`define Linv4 64'b1000000000100111101100101011100001011111000000010101001011101001
`define Linv5 64'b1000000000001000110110001101010101111010111010011100110110100011
`define Linv6 64'b1000000001111010001001110001011110110010100010011011100000110110
`define Linv7 64'b1000000011011000011110101100110100100111001010010001011100000100
`define Linv8 64'b1000000000100000000010000000001011011000001101101101010101011001
`define Linv9 64'b1000000011000000101000001111000010001000110011001010101011111111
`define Linv10 64'b1000000011011111110000000110100010100000010111001111000001110010
`define Linv11 64'b1000000000110010110111110011111111000000001010110110100011111000
`define Linv12 64'b1000000010100111001100101010110111011111111110010011111101001000
`define Linv13 64'b1000000011111010101001111100101000110010110000011010110101111111
`define Linv14 64'b1000000010001000010110001000010111111010000110111110111101111000
`define Linv15 64'b1000000010100000100010001010101001011000010011101000010111001000
`define Linv16 64'b1000000001011000111110101110111110100111010101101100101011110010
`define Linv17 64'b1000000010100010010111011101010010010101000110111001010011000100
`define Linv18 64'b1000000000101000110100000011100110100010110011001000101101101011
`define Linv19 64'b1000000010010101111011011011010000011111110000011011110001100001
`define Linv20 64'b1000000011101101000111111011110001100000111110010110010001110001
`define Linv21 64'b1000000001100000001010000001111011010000010111000011100110100110
`define Linv22 64'b1000000000011111011000000110010000101000001010110001111001110011
`define Linv23 64'b1000000001011101100101011001010011101101010101101011010010010110
`define Linv24 64'b1000000011010000101000101000101101011101010011101101010001111100
`define Linv25 64'b1000000010000010010101011001000101001101110100111101101111100101
`define Linv26 64'b1000000011010010011101111101000110010000101001001111101111111101
`define Linv27 64'b1000000001110111100100001111101110000010101111101111111000011101
`define Linv28 64'b1000000001010101010011011101101110010111001011101111011011000111
`define Linv29 64'b1000000001001101100101111111011000111000001100110100100100011010
`define Linv30 64'b1000000010010111001110000100100111010010100001101010000100001111
`define Linv31 64'b1000000000111000110100101010000101110111011000111101000101100010
`define Linv32 64'b1000000010010000100000101111111001010101101100011001000110110101
`define Linv33 64'b1000000001010010111101111111010000010000011001101001110011000110
`define Linv34 64'b1000000000000010110101011100011011001101100111000100001101100110
`define Linv35 64'b1000000011010101110011010100001100010111011011001010110011001011
`define Linv36 64'b1000000011110111000100001001110000000010110010110110110001000011
`define Linv37 64'b1000000000010000000000100110110011010101111101001100011010101100
`define Linv38 64'b1000000010111000010100101100101111110111101011001111010001101100
`define Linv39 64'b1000000000010111101110000110011001010010010000111100101110011100
`define Linv40 64'b1000000011001101000101111010110010111000110001100110011011110100
`define Linv41 64'b1000000010101000010100000100000100100010110001100111100111001111
`define Linv42 64'b1000000000100010110111011010101100010101101011001101110001110101
`define Linv43 64'b1000000001010000001000100111100111011101010000111010101111000010
`define Linv44 64'b1000000011011101000101011101110001101101011001100100110001000101
`define Linv45 64'b1000000001101101100111111100111011100000111101001001101101000010
`define Linv46 64'b1000000011100000101010001101011001010000011011000100000111000101
`define Linv47 64'b1000000010011111111000001001101110101000100111001101011011110101
`define Linv48 64'b1000000000010101011011010100110010011111110010111100111001001111
`define Linv49 64'b1000000000001111011000100010001011111101110011001101110101111011
`define Linv50 64'b1000000001100010111111011101110100011101010011100001010101111110
`define Linv51 64'b1000000011111101000111010001010110110101000110110110110100010001
`define Linv52 64'b1000000000011010000011110101000001100010010111000010001001010001
`define Linv53 64'b1000000000011101101101010110110111100101010101101001111101011011
`define Linv54 64'b1000000011000111000110101010100000001111001010110101000000100001
`define Linv55 64'b1000000010110101111001011001111111000111110000011110000001110110
`define Linv56 64'b1000000011100101110001111110000000011010111110011010100011001001
`define Linv57 64'b1000000010001111111000101100111101111101101111101100001001011000
`define Linv58 64'b1000000001111101100111010111010100110101110100110100010110100111
`define Linv59 64'b1000000011100010011111011100001010011101101100010111010111111010
`define Linv60 64'b1000000010011010100011111100010111100010101001001100111110001000
`define Linv61 64'b1000000001100101010001110100001010011010100001101111010111000000
`define Linv62 64'b1000000000110101011001010100111101000111001100110100001011011111
`define Linv63 64'b1000000001000111100110101111010110001111011000111100010110100000
`define Linv64 64'b1000000010011101001101010100010101100101001011100100111100110010
`define Linv65 64'b1000000001101010001001011010101101100111101001001101110010100010
`define Linv66 64'b1000000010010010010101111100111010011000110100111001101111101101
`define Linv67 64'b1000000001010111100110001001101101011010001011101101011000011111
`define Linv68 64'b1000000000100101011001111101110010010010101111100100110001011101
`define Linv69 64'b1000000001011010001011110100000101101010100001100111100100101000
`define Linv70 64'b1000000000101111011010100111100100100101011000111010101111010000
`define Linv71 64'b1000000001100111100100100100110001010111101100011100111010010101
`define Linv72 64'b1000000010011000010110101101011000101111001100110100000101100000
`define Linv73 64'b1000000000010010110101111000101100011000010110011101010010110110
`define Linv74 64'b1000000011101010101001010110010011100111001010010001111011011001
`define Linv75 64'b1000000011010111000110001101010011011010101000111001010001101001
`define Linv76 64'b1000000010100101111001110001111000010010100010010011100100100011
`define Linv77 64'b1000000011100111000100100011100111010111000000011000101110000100
`define Linv78 64'b1000000000011000110110101001010010101111000001001011010010101001
`define Linv79 64'b1000000011011010101011111011010011101010001101101011110000001001
`define Linv80 64'b1000000010101111111010101011110010100101111010010110010010000001
`define Linv81 64'b1000000011110010011111110100000101001000010000000111100111100111
`define Linv82 64'b1000000001001000111110001010101101110010000010001101110011010111
`define Linv83 64'b1000000011001000011110001001101111110010101100101101011011101010
`define Linv84 64'b1000000001110010111111110100110011001000011110101100111011011010
`define Linv85 64'b1000000011111000011100101101110011111111110110000100110000011000
`define Linv86 64'b1000000011111111110010001100111001111000001001111001101110101111
`define Linv87 64'b1000000001111111010010000111100111111000001000001010101100010010
`define Linv88 64'b1000000001111000111100101101011001111111010111110100000110100101
`define Linv89 64'b1000000000101010000001011011001101101111101000110000011001001101
`define Linv90 64'b1000000000101101101111110011111011101000001010010011000101110111
`define Linv91 64'b1000000000000101011011110000011001001010000001001110001110010111
`define Linv92 64'b1000000001110000001010101010111000000101010110011011001101010101
`define Linv93 64'b1000000011101000011100000101001100101010000000011010111010000010
`define Linv94 64'b1000000001001010001011010010010010111111111010010011111011010010
`define Linv95 64'b1000000010111111111010000011000101110000100010010101001110010000
`define Linv96 64'b1000000001101111010010101110001100101101001101100010010000111000
`define Linv97 64'b1000000010101010100001010001110011101111011001101110110010011011
`define Linv98 64'b1000000010101101001111110010110001101000011011001110011010101011
`define Linv99 64'b1000000010000101111011111110110011001010110010110100011011010110
`define Linv100 64'b1000000011110000101010100111010010000101101011000001110011001110
`define Linv101 64'b1000000000111111011010001110011011110000110001100100101111011100
`define Linv102 64'b1000000011101111110010100100011010101101111101001100001101000001
`define Linv103 64'b1000000011001010101011011100001100111111100111000010110001111001
`define Linv104 64'b1000000001101000111100000100101110101010010000110111010001001100
`define Linv105 64'b1000000011001111110000100011100101110101110011011000101111101111
`define Linv106 64'b1000000001001111010000101011010011110101111101111011110001101000
`define Linv107 64'b1000000001110101010001011101010001001111101110001001010010101101
`define Linv108 64'b1000000011110101110001010110010011001111000000100001111010101010
`define Linv109 64'b1000000011000101110011110001111011000010110101010011100110000101
`define Linv110 64'b1000000001000010111101011011110011000101000100000110010011110000
`define Linv111 64'b1000000011000010011101011000101101000101000101111101010011001010
`define Linv112 64'b1000000001000101010011111001010001000010010100101011010000111111
`define Linv113 64'b1000000001010100000101000011111000110100001010110011000111111100
`define Linv114 64'b1000000000001011010101000010010000010100111110010011111011101011
`define Linv115 64'b1000000000010100001101000011000100111100010111000101001101000100
`define Linv116 64'b1000000011100100100111101011001110111001000110110000011011110001
`define Linv117 64'b1000000010111001000010111110001101010100110000010010010000100110
`define Linv118 64'b1000000000111100111001001010111010011110010011101011001111100001
`define Linv119 64'b1000000000110100001111000101001111100100110011001010111000010110
`define Linv120 64'b1000000010011110101110010000011000001011010101101110001111110011
`define Linv121 64'b1000000001001100110011101010111010011011000101111011001110110100
`define Linv122 64'b1000000011011100010011000101001111001110110011011010111010010100
`define Linv123 64'b1000000010101011110111000011000101001100110101010101001111010100
`define Linv124 64'b1000000011001110100110111011001111010110101110000000011010111100
`define Linv125 64'b1000000001000001011110010010010010101011000100000011111000111001
`define Linv126 64'b1000000001111001101010110011111011011100000000100011000110001011
`define Linv127 64'b1000000010011011110101100000011001000001010100101110001101100100
`define Linv128 64'b1000000011010110010000011110001101111001111101110010010000011110
`define Linv129 64'b1000000011110011001001100100100111101011010000001010000100010011
`define Linv130 64'b1000000001000100000101101111111011100001011110101001000110011001
`define Linv131 64'b1000000000010110111000011001000111110001001001111101101100000011
`define Linv132 64'b1000000000100110111010111010000111111100001000001101000110001110
`define Linv133 64'b1000000011110001111100111111011000100110010111110100100101101110
`define Linv134 64'b1000000011101011111111001101000101000100000010001111101110111011
`define Linv135 64'b1000000011100001111100011101101111110011101100101111011010001100
`define Linv136 64'b1000000011111100010001001111101100010110110110001111111011011110
`define Linv137 64'b1000000011101001001010010110110010001001110100111100011010100100
`define Linv138 64'b1000000000110110111010011001110000101001101100010110110001100011
`define Linv139 64'b1000000001011001101000110110011000000100011000111100101100101110
`define Linv140 64'b1000000000101001100010011100011000000001001011100100001110111110
`define Linv141 64'b1000000000000100001101101111010011101001101111101001110010000110
`define Linv142 64'b1000000010001001000000010100001101011001001100111010110010110001
`define Linv143 64'b1000000000000001010110011010110010100011100001100110011011010011
`define Linv144 64'b1000000010100011000001001100101100110110101001001111010000110011
`define Linv145 64'b1000000011011011111101101110111101001001010100101100101010101000
`define Linv146 64'b1000000011111110100100011010101011011011000101111000010110011111
`define Linv147 64'b1000000011111011111111101111000010010001110011011010101001101101
`define Linv148 64'b1000000010100001110100010011111111111011000000100110100011011101
`define Linv149 64'b1000000011010001111110110110100011111110110101011111000000010101
`define Linv150 64'b1000000010010001110110111000010111110110101110001110111111100000
`define Linv151 64'b1000000001001001101000011010110111010001000100000011111100100010
`define Linv152 64'b1000000011110110010010011100101010100001111101111010110101010000
`define Linv153 64'b1000000011011110100110010110110100000011000001001001111101100101
`define Linv154 64'b1000000000010011100011100010001010111011000000011101110101111101
`define Linv155 64'b1000000010011001000000111001111110001100001101101110000001000111
`define Linv156 64'b1000000000000011100011001110000001101110111010011010100010011010
`define Linv157 64'b1000000010001110101110111101110111011110010110010001010110011101
`define Linv158 64'b1000000001101110000100110101000010001110100010010010001011100010
`define Linv159 64'b1000000010001100011011101010100000010011001010010101000010001111
`define Linv160 64'b1000000010111011110111100001010110011001101000110110110100110101
`define Linv161 64'b1000000010100100101111101101010110110001111110011100110100011011
`define Linv162 64'b1000000010000110011000110001000010100100010101100000001011001100
`define Linv163 64'b1000000000110011100001101111011101100011000110110001000001011100
`define Linv164 64'b1000000010111110101100011100110111010011001010110001011101010110
`define Linv165 64'b1000000011010011001011101011100000110011110011000101001011111001
`define Linv166 64'b1000000010110001110100110001011100101110010111001011100011000001
`define Linv167 64'b1000000000101110001100110101001010000110010011101111011100101011
`define Linv168 64'b1000000001100011101001000000001010111110110000011101010101001110
`define Linv169 64'b1000000001001011011101001010100000011100000000100101000010101110
`define Linv170 64'b1000000001000110110000110001010100101100101110000110110100100100
`define Linv171 64'b1000000000011100111011000010001001000110110011011101110100000110
`define Linv172 64'b1000000011000011001011000110110111100110010100101001111100111110
`define Linv173 64'b1000000011101100010001101101110111000011000101110001010111100011
`define Linv174 64'b1000000000101100111001101001111101001011111101111110000000110001
`define Linv175 64'b1000000011100110010010111110000001110100000100001010100001010011
`define Linv176 64'b1000000001110100000111000101000011101100110101010010001010110011
`define Linv177 64'b1000000001011110000110011010101010000011010110011000010101010111
`define Linv178 64'b1000000010010011000011100011111100111011001010010110100000100101
`define Linv179 64'b1000000000011001100000111000010100001100101000111110111110011000
`define Linv180 64'b1000000010000011000011001110111111101110000001001100101001011010
`define Linv181 64'b1000000000111011010111101111000000011001000000011010101010010010
`define Linv182 64'b1000000011101110100100111010110100001110111010010011111101101010
`define Linv183 64'b1000000000001100111011101100101010010011001101101010110100101111
`define Linv184 64'b1000000000001110001110110110100001011110100010011111000001100111
`define Linv185 64'b1000000001011011011101100100001011001001010000001111010100111011
`define Linv186 64'b1000000001111011011111100111010100010001001001110100010111101110
`define Linv187 64'b1000000001111110000100010100010101011011101100100100111110010011
`define Linv188 64'b1000000000100001010100011100111101111011110110001100001010000011
`define Linv189 64'b1000000001110110110010011111010100100001001000001100010101011110
`define Linv190 64'b1000000000010001010110110100111101110110010111110100001000001110
`define Linv191 64'b1000000011001001001000011100010101010001000010001100111100011001
`define Linv192 64'b1000000001010001011110111100001001111110011110100111010100001100
`define Linv193 64'b1000000011001011111101000001011110011100110101011011100011110111
`define Linv194 64'b1000000011000110010000110001000010101100010100100000001011001101
`define Linv195 64'b1000000011110100100111001011100001101100110011010101001000010000
`define Linv196 64'b1000000001100110110010111100110111110100000000100001011101010010
`define Linv197 64'b1000000010101100011001101101010111001011000100001100110110111000
`define Linv198 64'b1000000001000011101011000000001001100110111101111101010100010111
`define Linv199 64'b1000000001101100110001101111011101000011101110000001000011010101
`define Linv200 64'b1000000010011100011011000101001011000110000101111111011100000010
`define Linv201 64'b1000000000100100001111100100111100110001011011000100001011010001
`define Linv202 64'b1000000000000110111000110111010100100100111101000100010101001001
`define Linv203 64'b1000000010110011000001101100001011100011110010110111010111110110
`define Linv204 64'b1000000000111110001100010100001001010011110001101111010111111011
`define Linv205 64'b1000000011100011001001000100010100111110100111000100111110100001
`define Linv206 64'b1000000010101110101100111100111100000110011001101100001011011011
`define Linv207 64'b1000000001010011101011101100010110110011101011001100111110010001
`define Linv208 64'b1000000000110001010100111111010110101110010000111100010111111110
`define Linv209 64'b1000000001101001101010010010110000001001001100111110011000010100
`define Linv210 64'b1000000010110110011010011100001110101001001011100010110001010100
`define Linv211 64'b1000000010101001000010011110011010000001100001100100101100110100
`define Linv212 64'b1000000011011001001000110001110010000100101111101110110010011110
`define Linv213 64'b1000000000100011100001001110110010110110101100010100011010111001
`define Linv214 64'b1000000010000001110110010111010000100011101001000001110011100100
`define Linv215 64'b1000000000001001100000010100101111011001011000110111010000111100
`define Linv216 64'b1000000010000100101101100100011001101001110100111100001100001011
`define Linv217 64'b1000000011001100010011101010110000011011010000000110011000100111
`define Linv218 64'b1000000001011100110011000100001101001110010111111010110001111010
`define Linv219 64'b1000000000101011010111001100011011001100101100100100001111011000
`define Linv220 64'b1000000001001110000110110110011001010110001000001100101110110010
`define Linv221 64'b1000000001010110110000011111010011111001110110001001110001000000
`define Linv222 64'b1000000000011011010101101100101111000001000010001111010001011111
`define Linv223 64'b1000000011111001001010110110110001011100001001111100011000001000
`define Linv224 64'b1000000011000001111110011001110000101011011110100110110000100000
`define Linv225 64'b1000000010010110011000011110011001110001010000000100101111101000
`define Linv226 64'b1000000001110011101001100001110001101011110110001110110000000101
`define Linv227 64'b1000000011000100100101100010110001100001010111111110011010111111
`define Linv228 64'b1000000010100110011010111110110001111100011110100100011001101111
`define Linv229 64'b1000000001111100110001001100001110010110101100100010110000101101
`define Linv230 64'b1000000001100001011100010100101101110011001000000111010001110000
`define Linv231 64'b1000000001101011011111000100011011000100001001111100001101001010
`define Linv232 64'b1000000001110001011100110111010010100110000010000001110000101010
`define Linv233 64'b1000000011010100100101001111111010110100110010111001000100101100
`define Linv234 64'b1000000010001011110101001111101110010100011001101111111011000011
`define Linv235 64'b1000000010010100101101001001000110111100111101001101101111100110
`define Linv236 64'b1000000001100100000111100100100100111001110001101010000100011100
`define Linv237 64'b1000000000011110001110011010000110001011010000111101000111101100
`define Linv238 64'b1000000010110100101111001101101101100100100111001111011001001011
`define Linv239 64'b1000000010111100011001001111011000011110011011000100100101110100
`define Linv240 64'b1000000000111001100010111101000111010100101011001111101101000110
