`define w1 15'b110001100000000
`define w2 15'b100111101000000
`define w3 15'b101001000000000
`define w4 15'b111100000000000
`define w5 15'b100111011000000
`define w6 15'b111110001000000
`define w7 15'b100010111000000
`define w8 15'b110111011000000
`define w9 15'b111100010000000
`define w10 15'b111001001000000
`define w11 15'b101001100000000
`define w12 15'b111010100000000
`define w13 15'b110000100000000
`define w14 15'b100001100000000
`define w15 15'b110011101000000
`define w16 15'b110101100000000
`define w17 15'b110100001000000
`define w18 15'b111110111000000
`define w19 15'b111000101000000
`define w20 15'b110011100000000
`define w21 15'b110001010000000
`define w22 15'b100101001000000
`define w23 15'b101011100000000
`define w24 15'b110010101000000
`define w25 15'b110101110000000
`define w26 15'b110010001000000
`define w27 15'b101010100000000
`define w28 15'b110101100000000
`define w29 15'b110000111000000
`define w30 15'b101100010000000
