`define Linv1 64'b1000000001000000001000000001000000001000000001000000001000000001
`define Linv2 64'b1000000011000000101000001111000010001000110011001010101011111111
`define Linv3 64'b1000000010100010010111011101010010010101000110111001010011000100
`define Linv4 64'b1000000010000010010101011001000101001101110100111101101111100101
`define Linv5 64'b1000000001010010111101111111010000010000011001101001110011000110
`define Linv6 64'b1000000010101000010100000100000100100010110001100111100111001111
`define Linv7 64'b1000000000001111011000100010001011111101110011001101110101111011
`define Linv8 64'b1000000010001111111000101100111101111101101111101100001001011000
`define Linv9 64'b1000000001101010001001011010101101100111101001001101110010100010
`define Linv10 64'b1000000000010010110101111000101100011000010110011101010010110110
`define Linv11 64'b1000000011110010011111110100000101001000010000000111100111100111
`define Linv12 64'b1000000000101010000001011011001101101111101000110000011001001101
`define Linv13 64'b1000000010101010100001010001110011101111011001101110110010011011
`define Linv14 64'b1000000011001111110000100011100101110101110011011000101111101111
`define Linv15 64'b1000000001010100000101000011111000110100001010110011000111111100
`define Linv16 64'b1000000001001100110011101010111010011011000101111011001110110100
`define Linv17 64'b1000000011110011001001100100100111101011010000001010000100010011
`define Linv18 64'b1000000011101001001010010110110010001001110100111100011010100100
`define Linv19 64'b1000000011011011111101101110111101001001010100101100101010101000
`define Linv20 64'b1000000011011110100110010110110100000011000001001001111101100101
`define Linv21 64'b1000000010100100101111101101010110110001111110011100110100011011
`define Linv22 64'b1000000001001011011101001010100000011100000000100101000010101110
`define Linv23 64'b1000000001011110000110011010101010000011010110011000010101010111
`define Linv24 64'b1000000001011011011101100100001011001001010000001111010100111011
`define Linv25 64'b1000000011001011111101000001011110011100110101011011100011110111
`define Linv26 64'b1000000000100100001111100100111100110001011011000100001011010001
`define Linv27 64'b1000000001101001101010010010110000001001001100111110011000010100
`define Linv28 64'b1000000011001100010011101010110000011011010000000110011000100111
`define Linv29 64'b1000000010010110011000011110011001110001010000000100101111101000
`define Linv30 64'b1000000011010100100101001111111010110100110010111001000100101100
