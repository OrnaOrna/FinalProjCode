`define w1 16'b1100011000000000
`define w2 16'b1001111010000000
`define w3 16'b1010010000000000
`define w4 16'b1111000000000000
`define w5 16'b1001110110000000
`define w6 16'b1111100010000000
`define w7 16'b1000101110000000
`define w8 16'b1101110110000000
`define w9 16'b1111000100000000
`define w10 16'b1110010010000000
`define w11 16'b1010011000000000
`define w12 16'b1110101000000000
`define w13 16'b1100001000000000
`define w14 16'b1000011000000000
`define w15 16'b1100111010000000
`define w16 16'b1101011000000000
`define w17 16'b1101000010000000
`define w18 16'b1111101110000000
`define w19 16'b1110001010000000
`define w20 16'b1100111000000000
`define w21 16'b1100010100000000
`define w22 16'b1001010010000000
`define w23 16'b1010111000000000
`define w24 16'b1100101010000000
`define w25 16'b1101011100000000
`define w26 16'b1100100010000000
`define w27 16'b1010101000000000
`define w28 16'b1101011000000000
`define w29 16'b1100001110000000
`define w30 16'b1011000100000000
