`define W21_1 64'b0100011101011001010101101101000111111110011010010100111000110001
`define W21_2 64'b1000011101110001000010100011011110001101110100001111111001001101
`define W21_3 64'b0100101001101001110010111000110001111000001001001101100001000100
`define W21_4 64'b1010010000110011101100011011001011111011000010101000000110011011
`define W21_5 64'b0010011101001111001000010101000000011001010011011000000101101101
`define W21_6 64'b1110111001100100101000101011001011101100010101001010011101000111
`define W21_7 64'b0001011000011110001010100000100011010110101111111100111000111011
`define W21_8 64'b1011011110111001010110101011010111010110000101101010011000011001
`define W21_9 64'b0101011111100000111000011010000110010000111111000000100100011011
`define W21_10 64'b0101011101111111010110001000001101110111111110001001001110110101
`define W21_11 64'b0000000111100110010101001001111000001111001001010000101011110011
`define W21_12 64'b0110101000111111000110010110000000010001000101110110001110101110
`define W21_13 64'b1011001101101001100110101000101101001001010010111111011001000111
`define W21_14 64'b1110111010101111011011101001111110011011100011010110101100101100
`define W21_15 64'b1000111110010110000111101110110001111000110000001000000010110010
`define W21_16 64'b0111011011011111101010010110111001111110011010011110011001010010
`define W21_17 64'b0011101011111100101111111010111100011000011010001101001000111101
`define W21_18 64'b1001110111100100111111001111110100100001100000011010111100101110
`define W21_19 64'b1101000101000001110000001001100101101111111010011011111000001000
`define W21_20 64'b1010111010101100110111001100101010011001000010110000111011111011
`define W21_21 64'b1000011100001100000011100011110001001100000101111001011000010100
`define W21_22 64'b1010100101110001010001100101010101110011110000111101100010101111
`define W21_23 64'b1000010010101110101001101000001101010010001100111101110111011000
`define W21_24 64'b1111111010100001010101010001000101000110110100111111010110100110
`define W21_25 64'b0101110110110110100001000001100010101000000111101000000100001111
`define W21_26 64'b1100101101101010110010100010011011111000000011010001000001010100
`define W21_27 64'b0110011001001111011000000010001011000001101011010110110011110000
`define W21_28 64'b1010110011101010000101001101011100010101110011101010011001000111
`define W21_29 64'b1001111101011000100101110100110000100100110100000001000010110011
`define W21_30 64'b0100110010011110111010011011010100011111100001000001011011010110
