`define W21_1 40'b0101100001000110010010011100111011100001
`define W21_2 40'b1100101000111100010001110111101011000000
`define W21_3 40'b1000110110101110000011000100101110111111
`define W21_4 40'b0101000111000110010001000100011100001110
`define W21_5 40'b0100000000101000010001100011011101111110
`define W21_6 40'b1101101101010001100101111000011111011001
`define W21_7 40'b1010110010100100100100001011001001101100
`define W21_8 40'b1110011011101000000010111110010010000111
`define W21_9 40'b0010111010011001100110001101100011101001
`define W21_10 40'b0100000001101000010011111001010001100000
`define W21_11 40'b0011010111010010011000001010101000111011
`define W21_12 40'b1100010010010001101101111100111010111111
`define W21_13 40'b0001001111001001001110100010101111101001
`define W21_14 40'b0101110100011100110111010010110000101000
`define W21_15 40'b0100001001011011110100110010000110110101
`define W21_16 40'b0110011011001111101110010111111001101110
`define W21_17 40'b0111101110111101111111101110111001011001
`define W21_18 40'b1101011010101111101101111011011001101010
`define W21_19 40'b1000010100010101100101001100110100111011
`define W21_20 40'b0011111000111100010011000101101000001001
`define W21_21 40'b1101010101011110010111000110111000011110
`define W21_22 40'b0111011010101110100110011000101010101100
`define W21_23 40'b0100011001101100011001000100000110010000
`define W21_24 40'b1100001110011100011010000010110001111011
`define W21_25 40'b1110010100001110001111001010000000010000
`define W21_26 40'b1101110101111100110111000011000011101110
`define W21_27 40'b1110000111001000111001111010010101000110
`define W21_28 40'b0101110100011011111001010010011011100100
`define W21_29 40'b0100011110000000010011111001010011111100
`define W21_30 40'b0000101111011001101011101111001001011000
