`define w1 13'b1100011000000
`define w2 13'b1001111010000
`define w3 13'b1010010000000
`define w4 13'b1111000000000
`define w5 13'b1001110110000
`define w6 13'b1111100010000
`define w7 13'b1000101110000
`define w8 13'b1101110110000
`define w9 13'b1111000100000
`define w10 13'b1110010010000
`define w11 13'b1010011000000
`define w12 13'b1110101000000
`define w13 13'b1100001000000
`define w14 13'b1000011000000
`define w15 13'b1100111010000
`define w16 13'b1101011000000
`define w17 13'b1101000010000
`define w18 13'b1111101110000
`define w19 13'b1110001010000
`define w20 13'b1100111000000
`define w21 13'b1100010100000
`define w22 13'b1001010010000
`define w23 13'b1010111000000
`define w24 13'b1100101010000
`define w25 13'b1101011100000
`define w26 13'b1100100010000
`define w27 13'b1010101000000
`define w28 13'b1101011000000
`define w29 13'b1100001110000
`define w30 13'b1011000100000

