`define w1 12'b110001100000
`define w2 12'b100111101000
`define w3 12'b101001000000
`define w4 12'b111100000000
`define w5 12'b100111011000
`define w6 12'b111110001000
`define w7 12'b100010111000
`define w8 12'b110111011000
`define w9 12'b111100010000
`define w10 12'b111001001000
`define w11 12'b101001100000
`define w12 12'b111010100000
`define w13 12'b110000100000
`define w14 12'b100001100000
`define w15 12'b110011101000
`define w16 12'b110101100000
`define w17 12'b110100001000
`define w18 12'b111110111000
`define w19 12'b111000101000
`define w20 12'b110011100000
`define w21 12'b110001010000
`define w22 12'b100101001000
`define w23 12'b101011100000
`define w24 12'b110010101000
`define w25 12'b110101110000
`define w26 12'b110010001000
`define w27 12'b101010100000
`define w28 12'b110101100000
`define w29 12'b110000111000
`define w30 12'b101100010000
