`define w1 11'b11000110000
`define w2 11'b10011110100
`define w3 11'b10100100000
`define w4 11'b11110000000
`define w5 11'b10011101100
`define w6 11'b11111000100
`define w7 11'b10001011100
`define w8 11'b11011101100
`define w9 11'b11110001000
`define w10 11'b11100100100
`define w11 11'b10100110000
`define w12 11'b11101010000
`define w13 11'b11000010000
`define w14 11'b10000110000
`define w15 11'b11001110100
`define w16 11'b11010110000
`define w17 11'b11010000100
`define w18 11'b11111011100
`define w19 11'b11100010100
`define w20 11'b11001110000
`define w21 11'b11000101000
`define w22 11'b10010100100
`define w23 11'b10101110000
`define w24 11'b11001010100
`define w25 11'b11010111000
`define w26 11'b11001000100
`define w27 11'b10101010000
`define w28 11'b11010110000
`define w29 11'b11000011100
`define w30 11'b10110001000
