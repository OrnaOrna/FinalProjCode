interface multiplier_io;

endinterface