`define W21_1 48'b111010101111010011111011011111000101001111000100
`define W21_2 48'b001010111101110110100110100110110010000101111100
`define W21_3 48'b011010100100100111101011101011000101100000000100
`define W21_4 48'b110011010101101011011000110110111001001001100011
`define W21_5 48'b101100011101100110110111110001101000111111011011
`define W21_6 48'b011000011110101100101101001111010110001111011011
`define W21_7 48'b010101000101110001101000010010101001010011111101
`define W21_8 48'b000001000000101011101001000001100110010110100101
`define W21_9 48'b011000101101010111010100100101001010010111001001
`define W21_10 48'b001010110000001100100100111111110000101110000100
`define W21_11 48'b110110110011110010001110010001001101010111111111
`define W21_12 48'b111100101010011110000001111110001000100110001111
`define W21_13 48'b001100101110100000011011000010101100100011001010
`define W21_14 48'b101010011110100000101001110110001101110011001010
`define W21_15 48'b111111101110011101101111100111010000100110110001
`define W21_16 48'b001010111000001011110100001100110010001100110100
`define W21_17 48'b000101111101000110010010100000100011010101000101
`define W21_18 48'b111111111000011010011110100111110100001111100011
`define W21_19 48'b111101010110010111100100101111010100101111001101
`define W21_20 48'b111111101111110010001100100110101100100101011011
`define W21_21 48'b110010000100001101000001011100110000001101011000
`define W21_22 48'b110100100000101000111101001011100000100010111000
`define W21_23 48'b000111010011011100111111000110101100101110101010
`define W21_24 48'b011111010010001011010110100100101100010101010000
`define W21_25 48'b110101100011110100001111100100110010001110010101
`define W21_26 48'b010001101110011101000111101010110111010110000000
`define W21_27 48'b011111000101010101111010001110001101101110110111
`define W21_28 48'b100110001101111000100000111000110010000111111010
`define W21_29 48'b111001110010000011101111001101000101110010101000
`define W21_30 48'b000001101101010010100011111111110101010111001110
