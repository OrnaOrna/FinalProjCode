`define P 9'b100101101
`define Q 9'b110111101
`define PQ 17'b11000000000000001
`define d 8
`define W 256'b1001011000000000001001100000000000110110000000000110000000000000010101000000000011101110000000000111110100000000100011010000000001100101000000001000001000000000001100000000000011111010000000000110101100000000010000010000000001101110000000001001011100000000
`define w 16'b1010011000000000
`define pow1 256'b1000000000000000001000000000000000001000000000000000001000000000000000001000000000000000001000000000000000001000000000000000001011000000000000000011000000000000000011000000000000000011000000000000000011000000000000000011000000000000000011000000000000000011
`define pow2 256'b1000000000000000000010000000000000000000100000000000000000001000110000000000000000001100000000000000000011000000000000000000110010100000000000000000101000000000000000001010000000000000000010101111000000000000000011110000000000000000111100000000000000001111
`define pow4 256'b1000000000000000110000000000000010100000000000001111000000000000100010000000000011001100000000001010101000000000111111110000000010000000100000001100000011000000101000001010000011110000111100001000100010001000110011001100110010101010101010101111111111111111
`define r1 8'b11101111
`define r2 8'b11010110
`define r3 8'b01011001
`define r4 8'b10110101
`define r5 8'b11110000
`define r6 8'b01110010
`define r7 8'b00100010
`define L 64'b1000000000000100101100111010110100001100111110001101101000010100
`define L_inv 64'b1000000011110010011111110100000101001000010000000111100111100111
`define modPmat 64'b1001011001001011101100111100111111110001111011100111011110101101
`define mulL2 256'b0000010000000000000000100000000000000001000000000000000010000000000000000100000000000000001000000000000000010000000000000000100000000000000001000000000000000010000000000000000111000000000000000110000000000000001100000000000000011000000000000000110000000000
`define x_in 16'b0101011101010011
`define T2 16'b0001000100100101
`define t2 16'b1110011111101110
`define T3 16'b1010001111111110
`define t3 16'b0110101000000000
`define T12 16'b1100100001000000
`define t12 16'b1001100110010101
`define T14 16'b1110010010000101
`define T15 16'b1100011101010000
`define t14 16'b0100000011101100
`define t15 16'b0010110111100000
`define T240 16'b1111101111100000
`define t240 16'b1000010110001010
`define T254 16'b0011011111100111
`define t254 16'b0001000000011101
`define sbox_out 16'b1000000100000000
