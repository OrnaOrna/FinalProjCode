// Parameters used by the RAMBAM module with d=4 and P,Q chosen as per the original paper
`define P 9'b100101101
`define Q 9'b110111101
`define PQ 17'b11000000000000001
`define d 8
`define W 256'b1001011000000000001001100000000000110110000000000110000000000000010101000000000011101110000000000111110100000000100011010000000001100101000000001000001000000000001100000000000011111010000000000110101100000000010000010000000001101110000000001001011100000000
`define w 16'b1010011000000000
`define pow1 256'b1000000000000000001000000000000000001000000000000000001000000000000000001000000000000000001000000000000000001000000000000000001011000000000000000011000000000000000011000000000000000011000000000000000011000000000000000011000000000000000011000000000000000011
`define pow2 256'b1000000000000000000010000000000000000000100000000000000000001000110000000000000000001100000000000000000011000000000000000000110010100000000000000000101000000000000000001010000000000000000010101111000000000000000011110000000000000000111100000000000000001111
`define pow4 256'b1000000000000000110000000000000010100000000000001111000000000000100010000000000011001100000000001010101000000000111111110000000010000000100000001100000011000000101000001010000011110000111100001000100010001000110011001100110010101010101010101111111111111111
`define L 64'b1000000000000100101100111010110100001100111110001101101000010100
`define L_inv 64'b1000000011110010011111110100000101001000010000000111100111100111
`define modPmat 64'b1001011001001011101100111100111111110001111011100111011110101101
`define mulL2 256'b0000010000000000000000100000000000000001000000000000000010000000000000000100000000000000001000000000000000010000000000000000100000000000000001000000000000000010000000000000000111000000000000000110000000000000001100000000000000011000000000000000110000000000