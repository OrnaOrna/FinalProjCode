`define W11_1 64'b1111100001111100001111100001111110001111110001111110001111110001
`define W11_2 64'b1001100001001100001001100001001100001001000001000000001000000001
`define W11_3 64'b0101110011111100100111000010101010001001001001010110010110111101
`define W11_4 64'b1111001101010110001000001000101010001110001110001010010011100010
`define W11_5 64'b1001101010000000010110011100110110110010000001001011111100000101
`define W11_6 64'b0110000011110111000110001101110011111100101001111110101000110001
`define W11_7 64'b0111010111100101011001000000001001011100000001000001000010110000
`define W11_8 64'b1010001101110000000011110111011011010111110010001000101111101110
`define W11_9 64'b1000011001101101101101010010001100111011101001000001011000100000
`define W11_10 64'b0111000110011101011100001100110100111010001111000011000001000101
`define W11_11 64'b1001011000100110001101100110000001010100111011100111110110001101
`define W11_12 64'b0001001111010011101100001000001101011101010100010000101111001000
`define W11_13 64'b1010010101000000011101010100010100101110000001000010001100010100
`define W11_14 64'b1110100001001011110110110101011100100111101101101001111100100101
`define W11_15 64'b0011111110010110000101111001100000000111011011011111111000101011
`define W11_16 64'b0100000110000001000010010010010100100001010110101100001101101011
`define W11_17 64'b0000100111111100000101010101110101100111001100010111110010101100
`define W11_18 64'b0110111101001001111000000011101011100010000010000010100011111001
`define W11_19 64'b0011100101101011001101101011111100111100100000001100110100001000
`define W11_20 64'b0010010111011000001000000010110110111001111000000110001110110000
`define W11_21 64'b0110010101100001010000111111010111111011010110011011001111110010
`define W11_22 64'b0001001001010100100110010100010001001000010100001101000001100110
`define W11_23 64'b1001001110101011001100110001000000110100111011001010000110110010
`define W11_24 64'b0010011110011010000100010110110100110011000011101111111010001010
`define W11_25 64'b0101101010100110010111011010110100010010110111101010010101100011
`define W11_26 64'b0101001111001100110001100111101010011110010001101000111011001111
`define W11_27 64'b0111000111000110100100010101010000111011000001001111001111011001
`define W11_28 64'b0011111101000000010010001010010001100000000011010000001001000001
`define W11_29 64'b0010100101111011001010111011100101001010111001101010000001000011
`define W11_30 64'b0100000101010111001010001100011011011000000101010100111100000111
